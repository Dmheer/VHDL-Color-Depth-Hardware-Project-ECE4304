----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/06/2019 03:15:00 PM
-- Design Name: 
-- Module Name: PROM_IMG - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.math_real.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PROM_IMG is
    generic(DEPTH    :positive:= 450; 
            DATA_SIZE:positive:= 1600
           );
    Port   ( addr    : in  STD_LOGIC_VECTOR (integer(ceil(log2(real(449))))-1 downto 0);
             PROM_OP : out STD_LOGIC_VECTOR (1599 downto 0)
           );
end PROM_IMG;

architecture Behavioral of PROM_IMG is

type mem_type is array (0 to 449) of std_logic_vector (1599 downto 0);
signal mem: mem_type:= (
"1111110110101111111111101001111111110110101111111111111111111111111111111111111111111111111111011010111111111010011111110110101111111111111111111111111111111111111111111010111111111111010010111111111111111111111010011111111111111111111111111111111111111111111111011001111111111101101111111111110110111111111111111111111111111111111111111111111111111010011111111111111111111110101111111111111110011111111111111111111111111111111111111111111111111101001111111111010001111111111101101011111111111111111111111111111111111111111111111010111111110100011111110100011111111111111111111111111111111111111110101111111111010011111111111111111111111111111111010001111111110110011111111111100001111111111111111111111111111111111111111111111110101111111110100111111110100111111111111111111111111111111111111101100111111111111010111111111111111111111111111111111111111101100111111111111110101111111111100111111111111111111111111111111111111111111111111111111001111111110110111111111110101111111111111111111111111111111111111111110110011111111111111101100111111111111111111111111111111111111111111101100111111111111110101111111111111010111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111101001111111110110101111111101101011111111111111111111111111111111111111111111111111110110101111111100100111111101101011111111111111111111111111111111111111110101101111111111110110101111111111111111110110100111111111111111111111111111111111111111111111111010111111111111101011111111111110101111111111111111111111111111111111111111111111111110101111111111111111111101100111111111111111100111111111111111111111111111111111111111111111111111101011111111111010011111111111101011111111111111111111111111111111111111111111110100011111111110101111111110101111111111111111111111111111111111111110001111111111010001111111111111111111111111111111111001111111111100101111111111011011111111111111111111111111111111111111111111111110101111111101001111111110101111111111111111111111111111111111111101100111111111011010111111111111111111111111111111111111111101101111111111111110011111111101101111111111111111111111111111111111111111111111111111011011111111110101111111110110011111111111111111111111111111111111111111111010111111111111111110101111111111111111111111111111111111111111111110101111111111110110011111111111100001111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111010010111111101101011111111011010011111111111111111111111111111111111111111111111111111101001111111101001111111010010111111111111111111111111111111111111111101101011111111111110100111111111111111111101001011111111111111111111111111111111111111111111111110101111111111111010111111111111001011111111111111111111111111111111111111111111111101000111111111111111111111101011111111111111101011111111111111111111111111111111111111111111111111010001111111110100011111111111010001111111111111111111111111111111111111111111110110101111111110000111111110101111111111111111111111111111111111111110001111111111011010111111111111111111111111111111110010111111111110101111111111100001111111111111111111111111111111111111111111111110101111111110101111111110100111111111111111111111111111111111111101100111111111010001111111111111111111111111111111111111111110101111111111110110011111111101011111111111111111111111111111111111111111111111111111100111111111010111111111111010111111111111111111111111111111111111111111111001111111111111111010011111111111111111111111111111111111111111110110011111111111111010111111111101000111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111101100111111111011010011111111110100111111111111111111111111111111111111111111111111111111010011111111010011111111110101111111111111111111111111111111111111111111010111111111111101001111111111111111111110010111111111111111111111111111111111111111111111111011011111111110110011111111111011001111111111111111111111111111111111111111111111111101001111111111111111111111010111111111111111001111111111111111111111111111111111111111111111111111010011111111100101111111111111010111111111111111111111111111111111111111111111110101111111111000111111101000111111111111111111111111111111111111101000111111111110010111111111111111111111111111111111010111111111110101111111111011001111111111111111111111111111111111111111111111110011111111110100111111110101111111111111111111111111111111111111110101111111111011001111111111111111111111111111111111111111110011111111111110100111111111110011111111111111111111111111111111111111111111111111101100111111111011011111111011001111111111111111111111111111111111111111111101001111111111111011001111111111111111111111111111111111111111111011001111111111111011001111111111100101111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111011010011111111110100111111111011001111111111111111111111111111111111111111111111111111110100111111110100111111101101001111111111111111111111111111111111111110110101111111111111010011111111111111111110110101111111111111111111111111111111111111111111111011001111111111101100111111111110100011111111111111111111111111111111111111111111111111001111111111111111111110110011111111111110110111111111111111111111111111111111111111111111111111000011111111101000111111111110100011111111111111111111111111111111111111111111101000111111111100011111111100111111111111111111111111111111111111111101011111111111010111111111111111111111111111111111000111111111110101111111111010001111111111111111111111111111111111111111111111110101111111110001111111110101111111111111111111111111111111111111110101111111111011011111111111111111111111111111111111111110110011111111111111010111111110110111111111111111111111111111111111111111111111111111110101111111111011111111111011001111111111111111111111111111111111111111101100111111111111111011011111111111111111111111111111111111111111111101011111111111101000111111111111010011111111101100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111101100111111111100001111111111010011111111111111111111111111111111111111111111111111111011001111111100001111111011010011111111111111111111111111111111111111111101011111111111110100111111111111111111101001011111111111111111111111111111111111111111111110110011111111111101001111111111110100111111111111111111111111111111111111111111111110110011111111111111111111110101111111111111110101111111111111111111111111111111111111111111111111110101111111101101011111111111110101111111111111111111111111111111111111111111111101011111111010001111111101011111111111111111111111111111111111111101011111111110100011111111111111111111111111111111010011111111110001111111111011001111111111111111111111111111111111111111111111110101111111110101111111110101111111111111111111111111111111111111110100111111111010011111111111111111111111111111111111111110101111111111111111001111111110101111111111111111111111111111111111111111111111111110110011111111101101111111111000111111111111111111111111111111111111111111110101111111111111111100111111111111111111111111111111111111111111101100111111111111110101111111111010001111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111011010111111110110101111111101101011111111111111111111111111111111111111111111111111110110011111110100011111110110100111111111111111111111111111111111111111111001111111111111100001111111111111111111010001111111111111111111111111111111111111111111111101101111111111111010111111111111100111111111111111111111111111111111111111111111111110100111111111111111111101100111111111111101100111111111111111111111111111111111111111111111111110000111111111010001111111111110100111111111111111111111111111111111111111111111100001111111011010111111011001111111111111111111111111111111111111101001111111110100011111111111111111111111111111110100111111111101101111111111010010111111111111111111111111111111111111111111111110101111111110001111110100011111111111111111111111111111111111111110011111111111101011111111111111111111111111111111111111110110111111111111011001111111111001111111111111111111111111111111111111111111111111110110111111111110011111111101100111111111111111111111111111111111111111111110011111111111111101011111111111111111111111111111111111111111110110101111111111110110111111111111101011111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111110110011111111101101001111111011010011111111111111111111111111111111111111111111111111101100111111101001011111111101001111111111111111111111111111111111111110110101111111111111010011111111111111111110110011111111111111111111111111111111111111111111111011011111111111110101111111111011001111111111111111111111111111111111111111111111101001011111111111111111111101001111111111111100111111111111111111111111111111111111111111111111111101011111111110010111111111111001011111111111111111111111111111111111111111111010001111111111010111111110001111111111111111111111111111111111111010001111111111110101111111111111111111111111111110100011111111101000111111111111010111111111111111111111111111111111111111111111110101111111110101111111110101111111111111111111111111111111111111110011111111111101011111111111111111111111111111111111111111001111111111111011011111111111011111111111111111111111111111111111111111111111111111001111111110100111111111110011111111111111111111111111111111111111111111010011111111111110110111111111111111111111111111111111111111111110110111111111111111001111111111110001111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111101001111111111010101111111110100111111111111111111111111111111111111111111111111111011001111111011010111111111000011111111111111111111111111111111111111111101011111111111110000111111111111111111110000111111111111111111111111111111111111111111111110110111111111101100111111111110100011111111111111111111111111111111111111111111111011001111111111111111111111010111111111111111001111111111111111111111111111111111111111111111111010001111111110100111111111111010001111111111111111111111111111111111111111111111010111111110100011111110110111111111111111111111111111111111111011010111111111110101111111111111111111111111111110100011111111101000111111111111010111111111111111111111111111111111111111111111110011111111110101111110110011111111111111111111111111111111111110100011111111111000111111111111111111111111111111111111111111001111111111111101011111111011011111111111111111111111111111111111111111111111111011001111111111001111111110110011111111111111111111111111111111111111111011001111111111111111010111111111111111111111111111111111111111111011001111111111111101011111111110110011111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111010110011111111101000111111111010001111111111111111111111111111111111111111111111111110110101111110110101111111110100111111111111111111111111111111111111111010110111111111111100001111111111111111111010001111111111111111111111111111111111111111111111101011111111111011001111111111101100111111111111111111111111111111111111111111111111010011111111111111111110110011111111111110110111111111111111111111111111111111111111111111111011010111111110110101111111111011010111111111111111111111111111111111111111111111010111111110110011111110110011111111111111111111111111111111111111010111111111110101111111111111111111111111111111110101111111101101011111111111010111111111111111111111111111111111111111111111110101111111100101111111100011111111111111111111111111111111111110110011111111101100111111111111111111111111111111111111111011001111111111111100111111111101011111111111111111111111111111111111111111111111111100111111111111001111111110110111111111111111111111111111111111111111111010001111111111111011001111111111111111111111111111111111111111111101011111111111101100111111111011010111111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101000111111111011010011111110110101111111111111111111111111111111111111111111111111111100111111101101001111111101001111111111111111111111111111111111111111110101111111111111010011111111111111111011010111111111111111111111111111111111111111111111101100111111111111010111111111101101011111111111111111111111111111111111111111111111100101111111111111111111110101111111111111110011111111111111111111111111111111111111111111111110110011111111110101111111111111010111111111111111111111111111111111111111111110100011111111110101111110110011111111111111111111111111111111111111010011111111101000111111111111111111111111111111110101111111111000111111111111010111111111111111111111111111111111111111111111110011111111110101111110110011111111111111111111111111111111111110110011111111101000111111111111111111111111111111111111111011011111111111101100111111111100111111111111111111111111111111111111111111111111111100111111111011011111111011011111111111111111111111111111111111111111101100111111111111111101011111111111111111111111111111111111111111101101111111111110110011111111111101011111111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111011010011111110110100111111101100111111111111111111111111111111111111111111111111111111010111111010010011111111000011111111111111111111111111111111111111111100111111111111110000111111111111111111110100111111111111111111111111111111111111111111111011011111111111110101111111111111010111111111111111111111111111111111111111111111111100111111111111111111111101011111111111101100111111111111111111111111111111111111111111111110110101111111111001011111111110100011111111111111111111111111111111111111111111100101111111101000111111110101111111111111111111111111111111111110100011111111101100111111111111111111111111111111110101111111111101011111111111010011111111111111111111111111111111111111111111110101111111110001111110110011111111111111111111111111111111111111010111111111101101111111111111111111111111111111111111111011011111111111110101111111101101111111111111111111111111111111111111111111111111101101111111111100111111111011011111111111111111111111111111111111111111110100111111111111101101111111111111111111111111111111111111111110110011111111111111010111111111101000111111111111111111111000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111110100111111101100001111111111010011111111111111111111111111111111111111111111111111110100111111110100111111101000111111111111111111111111111111111111111011010111111111111100011111111111111111111101011111111111111111111111111111111111111111111110101011111111111100111111111110110011111111111111111111111111111111111111111111111011001111111111111111111011001111111111111011011111111111111111111111111111111111111111111111110101111111111101011111111111110101111111111111111111111111111111111111111111110100111111101101011111101101111111111111111111111111111111111110110011111111111001011111111111111111111111111111110100111111111101011111111110110111111111111111111111111111111111111111111111110011111110110101111110100011111111111111111111111111111111111111010011111111110101111111111111111111111111111111111111111101011111111111110011111111101101111111111111111111111111111111111111111111111111110101111111101100111111111101111111111111111111111111111111111111111110110011111111111111110011111111111111111111111111111111111111111111010111111111111011001111111110110011111111111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111101001111111111010011111111110100111111111111111111111111111111111111111111111111101101011111111100001111111010010111111111111111111111111111111111111111110101111111111111010011111111111111111011010111111111111111111111111111111111111111111111101011111111111011010111111111101100111111111111111111111111111111111111111111111111010111111111111111111111010111111111111111001111111111111111111111111111111111111111111111111001011111111111001111111111101000111111111111111111111111111111111111111111101000111111111101011111101100111111111111111111111111111111111111110101111111111101011111111111111111111111111111101000111111111100011111111110100011111111111111111111111111111111111111111111110011111111100101111110110011111111111111111111111111111111111111010111111111110101111111111111111111111111111111111111101100111111111111110011111111101011111111111111111111111111111111111111111111111110110011111111110011111111101101111111111111111111111111111111111111111111010011111111111111000111111111111111111111111111111111111111111011011111111111101100111111111111010111111111111111111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111110110101111111101101011111111011001111111111111111111111111111111111111111111111111110110111111111010011111110110101111111111111111111111111111111111111101101011111111111110100111111111111111110110101111111111111111111111111111111111111111111111100111111111110110011111111111101011111111111111111111111111111111111111111111110100011111111111111111110110011111111111110110111111111111111111111111111111111111111111111111011001111111111010111111111111101011111111111111111111111111111111111111111111101011111111010011111111011011111111111111111111111111111111111110100111111111100011111111111111111111111111111101000111111111011001111111110110011111111111111111111111111111111111111111111110101111111110101111110100111111111111111111111111111111111111110010111111111110101111111111111111111111111111111111111101101111111111110110011111110110111111111111111111111111111111111111111111111111110110111111110110011111111110011111111111111111111111111111111111111111011001111111111111011001111111111111111111111111111111111111111111101011111111111110011111111111101011111111111111111111111101100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111101101011111111011010111111110110011111111111111111111111111111111111111111111111111101100111111110000111111101001011111111111111111111111111111111111111111010111111111101101011111111111111111101100111111111111111111111111111111111111111111111110111111111111110101111111111111010111111111111111111111111111111111111111111111101000111111111111111111101100111111111111101011111111111111111111111111111111111111111111111110010111111110100011111111111101001111111111111111111111111111111111111111111100001111111010001111111011011111111111111111111111111111111111110000111111111011001111111111111111111111111111111000111111111010001111111110100011111111111111111111111111111111111111111111110011111110110101111110110011111111111111111111111111111111111111001111111110110011111111111111111111111111111111111111101101111111111111010111111111101111111111111111111111111111111111111111111111111111001111111110110111111110110011111111111111111111111111111111111111111101011111111111111101011111111111111111111111111111111111111111110101111111111110110011111111101100111111111111111111111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111010011111111110100111111101101001111111111111111111111111111111111111111111111111011001111111011001111111011010111111111111111111111111111111111111111110101111111111010010011111111111111111010001111111111111111111111111111111111111111111111101011111111111101011111111111110101111111111111111111111111111111111111111111111101011111111111111111111101011111111111101100111111111111111111111111111111111111111111111110100111111111110001111111111111010111111111111111111111111111111111111111111110001111111111010111111011001111111111111111111111111111111111101000111111111010001111111111111111111111111111111101011111111010001111111110110011111111111111111111111111111111111111111111101011111111110101111110110111111111111111111111111111111111111010001111111110100011111111111111111111111111111111111111110011111111111111010111111110101111111111111111111111111111111111111111111111111110111111111111001111111111010111111111111111111111111111111111111111101100111111111111101000111111111111111111111111111111111111111110110111111111111011001111111111100101111111111111111111111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111110101011111111101001111111111010011111111111111111111111111111111111111111111111110110011111111000011111110110101111111111111111111111111111111111111101101011111111111110101111111111111111110100011111111111111111111111111111111111111111111111111111111111111001111111111101100111111111111111111111111111111111111111111111010001111111111111111111011001111111111111010111111111111111111111111111111111111111111111110110101111111111000111111111111010011111111111111111111111111111111111111111111010011111110100011111110101111111111111111111111111111111111101101011111111111010111111111111111111111111111111101001111111011010111111111100011111111111111111111111111111111111111111111101011111110110101111111010011111111111111111111111111111111111011001111111110100111111111111111111111111111111111111111110011111111111011001111111110111111111111111111111111111111111111111111111111111100111111111110111111111011001111111111111111111111111111111111111111110100111111111111110011111111111111111111111111111111111111111111001111111111111100111111111111010011111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111010101010101111111111111111111111111111111111111110101010101010101010101010101111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111011010111111110110101111111101100111111111111111111111111111111111111111111111111101100111111101001011111101101001111111111111111111111111111111111111011001111111111101101011111111111111111101000111111111111111111111111111111111111111111111111111111111110110011111111111101011111111111111111111111111111111111111111111111000011111111111111111111010011111111111011001111111111111111111111111111111111111111111111101000111111111101011111111110110011111111111111111111111111111111111111111110100111111110110011111110110111111111111111111111111111111111111101001111111111010111111111111111111111111111111101011111111110010111111111110101111111111111111111111111111111111111111111110011111111110011111110110011111111111111111111111111111111111010001111111111010111111111111111111111111111111111111110110011111111111011001111111110111111111111111111111111111111111111111111111111111100111111111100111111111011011111111111111111111111111111111111111110110011111111111110100011111111111111111111111111111111111111111011011111111111101100111111111010001111111111111111111110101111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000001111111111111111111111111111111111111111111111111111111111111010000000111111111111111111111111111111111111111111111110110000000000000100111111111111111111111110101010101010000000000000000000000000000100101011111111111111111111111111111111111111111111111111111111111111100001001111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110110101111111101101001111111011001111111111111111111111111111111111111111111111111111010111111010010111111011010111111111111111111111111111111111111110110101111111111010010111111111111111111011001111111111111111111111111111111111111111111111111111111111101100111111111111010111111111111111111111111111111111111111111111110101111111111111111111110101111111111110110111111111111111111111111111111111111111111111101101011111111010001111111111110101111111111111111111111111111111111111111110100011111111110001111110101011111111111111111111111111111111111101001111111111000111111111111111111111111111111100011111111111010111111111110101111111111111111111111111111111111111111111101011111110110101111111010111111111111111111111111111111111111101011111111111000111111111111111111111111111111111111110101111111111111101011111111111111111111111111111111111111111111111111111111111101101111111101100111111111100111111111111111111111111111111111111111110110111111111111110001111111111111111111111111111111111111111101100111111111110110011111111111101011111111111111111111110101101010000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000111111111111111111010101010111111111111111111111111111111111000000000011111111111111111111111111111111111111111101100000000000000000000010111111111111111111010000000000000000000000000000000000000000000000001001111111111111111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111",
"0111111111111111111111111111111111111111111111111111111111101001111111111010011111110110101111111111111111111111111111111111111111111111110110011111110100100111110110100111111111111111111111111111111111111101100111111111110100101111111111111111111010011111111111111111111111111111111111111111111111111111111111101001111111111110011111111111111111111111111111111111111111111101101011111111111111111101101111111111111110011111111111111111111111111111111111111111111111101001111111111010111111111101100111111111111111111111111111111111111111111110101111111101000111111110011111111111111111111111111111111111010001111111110100011111111111111111111111111111011001111111111010111111111110101111111111111111111111111111111111111111111101011111111110101111111010011111111111111111111111111111111111101001111111111010111111111111111111111111111111111111110110111111111111100111111111111111111111111111111111111111111111111111111111111110101111111110101111111101101111111111111111111111111111111111111111011001111111111111011001111111111111111111111111111111111111111110011111111111111010111111111110001111111111111111111111111101000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111111111111111111111111111111111111111111111111111111100000000000000111111111111111101000000000011111111111111111111111111111111000000000010111111111111111111111111111111111111111000000000000000000000000000101111111111111100000000000000000000000000000000000000000000000000000000111111111111100101111111111111111111111111111111111111100000000000011111111111111111111111111111111111",
"1001111111111111111111111111111111111111111111111111111111110110101111111110101011111101101011111111111111111111111111111111111111111111111111101001111101101011111111101001111111111111111111111111111111111111111010111111111101001001111111111111111110000111111111111111111111111111111111111111111111111111111111111010111111111101100111111111111111111111111111111111111111111111010011111111111111111111101011111111111101101111111111111111111111111111111111111111111111111001111111110100011111111111101011111111111111111111111111111111111111111101000111111101100111111101011111111111111111111111111111111111011010111111110110011111111111111111111111111111010001111111111000111111111110101111111111111111111111111111111111111111111110011111110110011111111010111111111111111111111111111111111111101011111111111010111111111111111111111111111111111111111001111111111101100111111111111111111111111111111111111111111111111111111111110110011111111110011111111110011111111111111111111111111111111111111111101011111111111111000111111111111111111111111111111111111111111010111111111111011011111111110110011111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111110100000000000000101111111111111100000000000010111111111111111111111111111111000000000000111111111111111111111111111111111110100000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000101111111110000000011111111111111111111111111111111111100000000000011111111111111111111111111111111111",
"1010101111111111111111111111111111111111111111111111111111111101101001111111011010111111111010011111111111111111111111111111111111111111111111111010111111011010011111111000111111111111111111111111111111111111110110101111111111010010111111111111111111100001111111111111111111111111111111111111111111111111111111110110011111111111011011111111111111111111111111111111111111111111111010111111111111111111111001111111111111010111111111111111111111111111111111111111111111111010011111111110101111111111011001111111111111111111111111111111111111111111000111111111101011111101100111111111111111111111111111111111111010111111111110101111111111111111111111111111110001111111111010111111111110101111111111111111111111111111111111111111111101011111111100011111111010111111111111111111111111111111111111101011111111010001111111111111111111111111111111111111011011111111111101100111111111111111111111111111111111111111111111111111111111110110111111111101111111110110011111111111111111111111111111111111111101100111111111111101101111111111111111111111111111111111111111011001111111111101101011111111011010111111111111111111111111111111010000000011111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000011111111111111111111111111111111111111111111111010000000000000000001111111111111110000000000000111111111111111111111111111111000000000010111111111111111111111111111111111000000000000000000000000000000000101111111111011000000000000000000000000000000000000000000000000000000000001011110100000000101111111111111111111111111111110100000000000000011111111111111111111111111111111111",
"1101101001111111111111111111111111111111111111111111111111111111011010011111110110100111111110100111111111111111111111111111111111111111111111111110100111110110100111111110100111111111111111111111111111111111111101101011111111110110011111111111111111111000111111111111111111111111111111111111111111111111111111111101100111111111110110111111111111111111111111111111111111111111111110101111111111111111110110011111111111111001111111111111111111111111111111111111111111111100101111111101000111111111110010111111111111111111111111111111111111111111101011111111100001111111100111111111111111111111111111111111111000011111111110101111111111111111111111111111110001111111110100011111111101101111111111111111111111111111111111111111111101011111110110101111111010111111111111111111111111111111111111100111111111011001111111111111111111111111111111111111111011111111111101101111111111111111111111111111111111111111111111111111111111111010111111110111111111111001111111111111111111111111111111111111111110101111111111110100011111111111111111111111111111111111111111101011111111111101101111111111101011111111111111111111111111111111100000001011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111101000000000000000000001111111111111100000000000000111111111111111111111111111111000000000011111111111111111111111111111111100000000000000000101010000000000000111111111111010000000000000000000000001010101010101010000000000000000000000011110100000000000111111111111111111111111111110100000000000000111111111111111111111111111111111111",
"1111011010111111111111111111111111111111111111111111111111111111111110000111111101101001111111011010111111111111111111111111111111111111111111111111011001111111100011111111101001111111111111111111111111111111111111011001111111111110100111111111111111110110101111111111111111111111111111111111111111111111111111111111010001111111111110011111111111111111111111111111111111111111111101100111111111111111111110101111111111110101111111111111111111111111111111111111111111111101001111111101101011111111110110011111111111111111111111111111111111111111010001111111111010111111010111111111111111111111111111111111110110011111111110001111111111111111111111111111111010111111110100011111111101100111111111111111111111111111111111111111111101011111110100011111111010111111111111111111111111111111111101100111111111010011111111111111111111111111111111111111011011111111111110101111111111111111111111111111111111111111111111111111111111011001111111111001111111111001111111111111111111111111111111111111110110011111111111110110111111111111111111111111111111111111111101101111111111110110111111111101000111111111111111111111111111111111010000001011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111100000000000000000000001111111111111110000000000000101111111111111111111111111111000000000011111111111111111111111111111110000000000000001001111111100000000000111111111111010000000000000010101010010111111111111111011010101000000000000011110100000000000001111111111111111111111111110000000000001011111111111111111111111111111111111111",
"1111111101100111111111111111111111111111111111111111111111111111111111011010011111110110011111110110011111111111111111111111111111111111111111111111110110011111011010011111111010011111111111111111111111111111111111110110101111111111011001111111111111111101101001111111111111111111111111111111111111111111111111111111110110111111111111100111111111111111111111111111111111111111111101101011111111111111111101100111111111111101111111111111111111111111111111111111111111111111101011111111101001111111111110011111111111111111111111111111111111111111111010111111111010111111010111111111111111111111111111111111111100011111111101100111111111111111111111111111111010111111110110011111111101100111111111111111111111111111111111111111111101111111110110011111111010111111111111111111111111111111111101100111111111101011111111111111111111111111111111111111100111111111110110011111111111111111111111111111111111111111111111111111111111011011111111010111111111101011111111111111111111111111111111111111111010111111111111011001111111111111111111111111111111111111111110011111111111011010111111110110011111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111110100000000000000000000001111111111111100000000000000000111111111111111111111111111000000000011111111111111111111111111111000000000000000011111111111100000000000011111111111100000000000000001111111111111111111111111111111111101100000000011110100000000000010111111111111111111111111000000000000001011111111111111111111111111111111111111",
"1011111111011001011111111111111111111111111111111111111111111111111111110110101111111101001011111111100101111111111111111111111111111111111111111111111101100111111110000111111101100111111111111111111111111111111111111101011011111111111010011111111111111111011010111111111111111111111111111111111111111111111111111111110110101111111111011011111111111111111111111111111111111111111111011010111111111111111111011001111111111111111111111111111111111111111111111111111111111111011001111111110010111111111110101111111111111111111111111111111111111111111000111111111000011111110111111111111111111111111111111111111110101111111111000111111111111111111111111111111010011111110100101111111101100111111111111111111111111111111111111111111111111111110110011111011010111111111111111111111111111111111101100111111111101011111111111111111111111111111111111111101111111111110110011111111111111111111111111111111111111111111111111111111111100111111111100111111111100111111111111111111111111111111111111111011001111111111111101001111111111111111111111111111111111111110110111111111111101011111111111010111111111111111111111111111111111101000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000101111111111111111111111111111111111100000000000000000000000001011111111111110000000000000001011111111111111111111111111000000000011111111111111111111111111100000000000000001111111111111000000000010111111111111110101000000001001111111111111111111111111111111111111110000000011111110000000000000011111111111111111111101000000000000001111111111111111111111111111111111111111",
"1010011111111101100111111111111111111111111111111111111111111111111111111101101001111111011010111111111010011111111111111111111111111111111111111111111111011001111111010001111111010001111111111111111111111111111111111111011001111111111110100111111111111111110100101111111111111111111111111111111111111111111111111111111111100111111111110101011111111111111111111111111111111111111111110110011111111111111111111010111111111111111111111111111111111111111111111111111111111111110010111111111010011111111101100111111111111111111111111111111111111111110110011111111100011111111111111111111111111111111111111111111110100111111111101011111111111111111111111111110100111111111110101111111101100111111111111111111111111111111111111111111111111111110110011111111010111111111111111111111111111111111110100111111111101011111111111111111111111111111111111101011111111111111010111111111111111111111111111111111111111111111111111111111110101111111101100111111101101111111111111111111111111111111111111111101011111111111101100111111111111111111111111111111111111111011001111111111101101111111111101001111111111111111111111111111111110110000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111100000000000000000000000000011111111111110000000000000000011111111111111111111111111000000000011111111111111111111111110000000000000000111111111111111100000000011111111111111111111100000000111111111111111111111111111111111111111110000000011111111100000000000011111111111111111111100000000000010111111111111111111111111111111111111111111",
"0110000111111111011010011111111111111111111111111111111111111111111111111111111010011111110110100111111101100111111111111111111111111111111111111111111111110110011111010100101111110100011111111111111111111111111111111111111110011111111111101001111111111111111101101011111111111111111111111111111111111111111111111111111111011001111111111101011111111111111111111111111111111111111111111110101111111111111111110110011111111111111111111111111111111111111111111111111111111111110100011111111110101111111111100111111111111111111111111111111111111111111110101111111110101111111111111111111111111111111111111111111101100111111111101011111111111111111111111111110100111111111110101111111111101111111111111111111111111111111111111111111111111111110100011111111010111111111111111111111111111111111110101111111111000111111111111111111111111111111111111101011111111111111010111111111111111111111111111111111111111111111111111111111110011111111101011111111110011111111111111111111111111111111111111101100111111111111110101111111111111111111111111111111111111111010111111111111110011111111101100111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111110000000000000000101000000000011111111111000000000000000000000111111111111111111111111000000000011111111111111111111111100000000000000011111111111111111010100000111111111111111111111100000000111111111111111111111111111111111111111100000000011111111010000000000000111111111111111110000000000000010111111111111111111111111111111111111111111",
"1101101010111111110110100111111111111111111111111111111111111111111111111111111101101011111111011001111111011001111111111111111111111111111111111111111111111101101011111101101011111101101011111111111111111111111111111111111101101011111111111010011111111111111111011001111111111111111111111111111111111111111111111111111111110110011111111101010111111111111111111111111111111111111111111101100111111111111111111110101111111111111111111111111111111111111111111111111111111111110110101111111110100111111111011011111111111111111111111111111111111111111110101111111101001111111111111111111111111111111111111111111111100111111111010011111111111111111111111111111100011111111110101111111111010111111111111111111111111111111111111111111111111111110110011111111001111111111111111111111111111111111110100111111101100111111111111111111111111111111111111101011111111111011001111111111111111111111111111111111111111111111111111111110110011111110110111111110110111111111111111111111111111111111111111110101111111111110110011111111111111111111111111111111111111101010111111111111010111111111110101111111111111111111111111111111111011000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111000000000011111111111000000000000000000000111111111111111111111111000000000011111111111111111111111000000000000001111111111111111111111111011111111111111111111111100000000111111111111111111111111111111111111110000000000011111111011000000000000111111111111111010000000000001001111111111111111111111111111111111111111111",
"1111110110100111111111101010111111111111111111111111111111111111111111111111111111011010011111110110101111110110010111111111111111111111111111111111111111111111111010111111010001111111011001111111111111111111111111111111111111011001111111111110101111111111111111110110011111111111111111111111111111111111111111111111111111111110101111111111110111111111111111111111111111111111111111111111011001111111111111111101101011111111111111111111111111111111111111111111111111111111111101000111111101101011111111111001111111111111111111111111111111111111111101000111111101101011111111111111111111111111111111111111111111100111111111011001111111111111111111111111111110101111111110001111111111100111111111111111111111111111111111111111111111111111110100011111011010111111111111111111111111111111111110101111111101001111111111111111111111111111111111111110011111111111011001111111111111111111111111111111111111111111111111111111110110111111110110111111110101111111111111111111111111111111111111110110111111111111011010111111111111111111111111111111111111110110011111111111011001111111110100111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111000000000000001111111000000000011111111111000000000000000000000001111111111111111111111000000000011111111111111111111100000000000000111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111000000000000111111111111110000000000001111111111111000000000000001111111111111111111111111111111111111111111111",
"1111111101011001111111110110101111111111111111111111111111111111111111111111111111111110100111111101001001111111101011111111111111111111111111111111111111111111111110101111110100010111110110011111111111111111111111111111111111111110101111111111101001111111111111111110000111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111010111111111111111111011001111111111111111111111111111111111111111111111111111111111111101011111111101001111111110110111111111111111111111111111111111111111111101011111111101011111111111111111111111111111111111111111111101011111111110001111111111111111111111111111100011111111110101111111111100111111111111111111111111111111111111111111111111111110110011111111001111111111111111111111111111111111100101111111110101111111111111111111111111111111111111101111111111111101011111111111111111111111111111111111111111111111111111111111001111111011001111111011001111111111111111111111111111111111111111010111111111111011011111111111111111111111111111111111111110110111111111111100111111111011001111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111000000000000001111111010000000010111111111000000000000000000000001111111111111111111111000000000011111111111111111110000000000000011111111111111111111111111111111111111111111111111111100000001011111111111111111111111111111111100000000000001111111111111111100000000000011111111101000000000000101111111111111111111111111111111111111111111111",
"1111111111110110011111111111101001011111111111111111111111111111111111111111111111111111100010111111111010011111110110011111111111111111111111111111111111111111111111011001111101101011111111101011111111111111111111111111111111111101101011111111111010011111111111111111101001111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111110110011111111111111111111010111111111111111111111111111111111111111111111111111111111111101001111111010001111111111110011111111111111111111111111111111111111111100001111111010001111111111111111111111111111111111111111111011011111111111010111111111111111111111111111110101111111101000111111111010111111111111111111111111111111111111111111111111111110100011111111001111111111111111111111111111111110110011111111110101111111111111111111111111111111111110101111111111111101011111111111111111111111111111111111111111111111111111111011011111111011001111111011011111111111111111111111111111111111111011011111111111101101011111111111111111111111111111111111111011001111111111110101111111111101011111111111111111111111111111111110100100000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111100000000000000111111111110000000000111111111100000000000000000000000011111111111111111111000000000011111111111111111100000000000001111111111111111111111111111111111111000000011111111111100000000111111111111111111111111111111110000000000000011111111111111111100000000000000111111100000000000000111111111111111111111111111111111111111111111111",
"1111111111111101101001111111111010101111111111111111111111111111111111111111111111111111110110101111111110100111111101100111111111111111111111111111111111111111111111110110111111011010011111011010111111111111111111111111111111111111111001111111111110101111111111111111111010111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111101100111111111111111110110011111111111111111111111111111111111111111111111111111111111110010111111111010011111111101011111111111111111111111111111111111111111111010111111011010111111111111111111111111111111111111111111111001111111111010111111111111111111111111111101101111111101100111111111010111111111111111111111111111111111111111111111111111110110011111111001111111111111111111111111111111110110011111111110011111111111111111111111111111111111110101111111111101100111111111111111111111111111111111111111111111111111111111101011111111101011111111100111111111111111111111111111111111111111101011111111111101101111111111111111111111111111111111111101100111111111110110011111111110101111111111111111111111111111111111110010010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000111111111010000000000111111111110000000000000000000000011111111111111111111000000000011111111111111111000000000000011111111111111111111110111010000000000000000001111111111100000000111111111111111111111111111011000000000000000111111111111111111111000000000000111110100000000000010111111111111111111111111111111111111111111111111",
"1111111111111111111000010111111101101001111111111111111111111111111111111111111111111111111111101001111111011001111111011001111111111111111111111111111111111111111111111101100111110110100111111110101111111111111111111111111111111111110110101111111111101011111111111111111110100111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111101011111111111111111101100111111111111111111111111111111111111111111111111111111111110100111111110100011111111111100111111111111111111111111111111111111111111010111111111010111111111111111111111111111111111111111111110101111111110110111111111111111111111111111101001111111101001011111111010111111111111111111111111111111111111111111111111111110100111111011001111111111111111111111111111111110110011111111100011111111111111111111111111111111111110111111111111101100111111111111111111111111111111111111111111111111111111101100111111101100111111101101111111111111111111111111111111111111101101111111111110110011111111111111111111111111111111111111101100111111111111001111111110110011111111111111111111111111111111111101001100000100111111111111111111111111111111111111111011101011101011101010101110101011101011101011101111111111111111111111111111111111111111111111111100000000000011111111111110000000010111111111100000000000000000000000000111111111111111111000000000011111111111111110000000000001111111111111101110110000000000000000000000000001111111111100000000111111111111111111111111110000000000000000011111111111111111111111110000000000001110000000000001011111111111111111111111111111111111111111111111111",
"1111111111111111111101101011111111111010011111111111111111111111111111111111111111111111111111111010101111110110101111111110011111111111111111111111111111111111111111111111011001111111101001111111101011111111111111111111111111111111111101101011111111111010111111111111111111101011111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111011001111111111111111111101011111111111111111111111111111111111111111111111111111111111110101111111110101111111111010111111111111111111111111111111111111111110100011111110100011111111111111111111111111111111111111111110101111111110100011111111111111111111111111101100111111111101011111111010101111111111111111111111111111111111111111111111111110100011111011001111111111111111111111111111111110110011111110100011111111111111111111111111111111111110111111111111110101111111111111111111111111111111111111111111111111111111101101111111110101111111110011111111111111111111111111111111111111110101111111111111010110111111111111111111111111111111111110110011111111111100111111111111010111111111111111111111111111111111110001111100000101111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111101000000000001111111111111110000000000111111111110000000000000000000000000111111111111111111000000000011111111111111100000000000011111111111111000000000000000000000000000000000000011111111100000001011111111111111111111011000000000000000000111111111111111111111111111000000000000010000000000001111111111111111111111111111111111111111111111111111",
"1111111111111111111111011010011111111101101011111111111111111111111111111111111111111111111111111101001011111101101001111111011011111111111111111111111111111111111111111111110110011111011010011111011010011111111111111111111111111111111111111010111111111110101111111111111111011010111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111110110011111111111111111011001111111111111111111111111111111111111111111111111111111111110100111111101101011111111111011111111111111111111111111111111111111110110101111110110101111111111111111111111111111111111111111110110111111111110101111111111111111111111111111000111111111001011111111010111111111111111111111111111111111111111111111111111110110111111011001111111111111111111111111111111111010011111110110011111111111111111111111111111111111010111111111111101101111111111111111111111111111111111111111111111111111111110011111111110101111111110111111111111111111111111111111111111111110111111111111011001111111111111111111111111111111111111111001111111111101101111111111101011111111111111111111111111111111110100011110000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111110000000000001111111111111110100000000001111111100000000110000000000000000001111111111111111000000000011111111111101100000000000111111111111010000000000000000000000000000000000000011111101100000000111111111111111110110000000000000000000111111111111111111111111111111100000000000000000000000101111111111111111111111111111111111111111111111111111",
"1111111111111111111111111101100101111111011010011111111111111111111111111111111111111111111111111111011010011111111010011111110101111111111111111111111111111111111111111111111101100111111110001111111110100111111111111111111111111111111111110101101111111111101011111111111111111110101111111111111111111111111111111111111111111111111111110100011111111111111111111111111111111111111111111111111111111110101111111111111111111010011111111111111111111111111111111111111111111111111111111111001011111111101011111111111001111111111111111111111111111111111111111110101111111110101111111111111111111111111111111111111111110101011111111110101111111111111111111111111111100111111101101011111111110111111111111111111111111111111111111111111111111111111000111111011001111111111111111111111111111111111010111111110100011111111111111111111111111111111111010111111111110110011111111111111111111111111111111111111111111111111111110110111111110110111111110101111111111111111111111111111111111111110111111111111111101011111111111111111111111111111111111111011011111111111110011111111101100111111111111111111111111111111111011010110100000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110100000000000111111111111111111100000000101111111110000000111100000000000000001011111111111111000000000011111111111110000000000011111111111111010000000000000000000000000000000000001011111110000000000111111111111101100000000000000000000011111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111011001011111111110101001111111111111111111111111111111111111111111111111110110100111111101101011111111111111111111111111111111111111111111111111111111111001011111101001111111101011111111111111111111111111111111111101100111111111011010111111111111111101101011111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111101100111111111111111111110101111111111111111111111111111111111111111111111111111111111011001111111010001111111110101011111111111111111111111111111111111111101100111111101000111111111111111111111111111111111111111111101011111111101101111111111111111111111111111101011111111101011111111110111111111111111111111111111111111111111111111111111110110011111011001111111111111111111111111111111111010111111111010111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111010111111110110111111011001111111111111111111111111111111111111010111111111111101000111111111111111111111111111111111111101010111111111110110111111110110011111111111111111111111111111111101101011110100001011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000101111111111111111110100000000001111111100000001111110000000000000000001111111111111000000000011111111111110000000000001111111111111010000000000000000000000000000000010101111111110000000000111111101101000000000000000000000000111111111111111111111111111111111111100000000000000000010111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101101011111111011010111111111111111111111111111111111111111111111111111111101001111111011010111111111111111111111111111111111111111111111111111111111110101111111000011111110110011111111111111111111111111111111111111010111111110110101111111111111111011010111111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111011001111111111111111101100111111111111111111111111111111111111111111111111111111111011001111111111010111111111101011111111111111111111111111111111111111111101011111101101011111111111111111111111111111111111111111101011111111101100111111111111111111111111111101011111111010001111111111111111111111111111111111111111111111111111111111111110100111111011001111111111111111111111111111111111010111111111010111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111001111111110111111111011011111111111111111111111111111111111111010111111111111110101111111111111111111111111111111111111101101111111111011011111111110110111111111111111111111111111111111101100111011000001011111111111111111111111111111111111111111111111010101000101000000000000000000000000010101000101010111111111111111111111111111111111111010000000000011111111111111111111100000000101111111110000001111111100000000000000000111111111111000000000011111111111110000000000111111111111111111100000000001010001000000000001111111111111110000000001010100100000000000000000000000000111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111011010011111110101101011111111111111111111111111111111111111111111111111110110101111110110100111111111111111111111111111111111111111111111111111111101011011111101000111111101100111111111111111111111111111111111110110011111111111101011111111111111110100011111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111010111111111111111111101011111111111111111111111111111111111111111111111111111111111000011111110100011111111101111111111111111111111111111111111111111111100011111111101011111111111111111111111111111111111111111111111111111111000111111111111111111111111111011011111111011001111111111111111111111111111111111111111111111111111111111111111010111111011001111111111111111111111111111111111001111111110010111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111011001111111011011111111100111111111111111111111111111111111111101101111111111110100111111111111111111111111111111111111110110111111111111100111111111011001111111111111111111111111111111110100011111100000001111111111111111111111111111111111111111111111111111111111111111101010101010101010101111111111111111111111111111111111111111111111111111100000000010111111110110101010101000000000101111111110000001111111111000000000000000000111111111000000000011111111110110000000000111111111111111111111101010011111110100000000001111111111111110000000000000000000000000000000000000001001111111111111111111111111111111111111111111100000000000001011111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111110101011111101011010111111111111111111111111111111111111111111111111111101101001111111011001111111111111111111111111111111111111111111111111111111111010011111010010111111101001111111111111111111111111111111111111100111111111011010111111111111111101101011111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111110011111111111111111011001111111111111111111111111111111111111111111111111111111111110101111111110101111111111111111111111111111111111111111111111111111011001111111101001111111111111111111111111111111111111111111111111111111100111111111111111111111111111011011111111010001111111111111111111111111111111111111111111111111111111111111111010111111011011111111111111111111111111111111011010111111111001111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111101011111111100111111101011111111111111111111111111111111111111110101111111111111001111111111111111111111111111111111111111001111111111110100111111111100111111111111111111111111111111111011010111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000101010100000000000000000000000000111111100000001111111111100000000000000000111111111000000000011111111111000000000001111111111111111111111111111111111110000000000101111111111111110000000000000000000000000000000000000011111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111011010011111110110100111111111111111111111111111111111111111111111111111111000011111110110101111111111111111111111111111111111111111111111111111111101100111110110101111110110011111111111111111111111111111111111010101111111110110101111111111111111011001111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111101100111111111111111110110011111111111111111111111111111111111111111111111111111111110000111111101000111111111111111111111111111111111111111111111111111111010111111110001111111111111111111111111111111111111111111111111111111101011111111111111111111111111010001111111011001111111111111111111111111111111111111111111111111111111111111111010111111010101111111111111111111111111111111011001111111010001111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111101100111111101010111111101011111111111111111111111111111111111110110011111111111010011111111111111111111111111111111111111011011111111110110011111111110011111111111111111111111111111111111101011110100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001001111110000001111111111110000000000000000001111111000000000011111111111000000000011111111111111111111111111111111111100000000000111111111111111110000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000101111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111110101101011111111101001111111111111111111111111111111111111111111111111111101101011111101101011111111111111111111111111111111111111111111111111111111011001111101001001111101100111111111111111111111111111111111110110011111111101101011111111111111111010011111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111101011111111111111111110101111111111111111111111111111111111111111111111111111111101101011111101100111111111111111111111111111111111111111111111111111111010011111111010111111111111111111111111111111111111111111111111111111011011111111111111111111111111111001111111010010111111111111111111111111111111111111111111111111111111111111111010111111011011111111111111111111111111111111011001111111011001111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111101101111111101011111111110011111111111111111111111111111111111111010111111111111000111111111111111111111111111111111111101100111111111011001111111110110111111111111111111111111111111111110100111010000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101000101111111111111100000000000000000000000000000000000000000000001011111100000001111111111111100000000000000000011111000000000011111111111000000000011111111111111111111111111111111101000000000010111111111111111101000000000000000000000000000000000000000111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111101010111111110110100111111111111111111111111111111111111111111111111111011010011111111010011111111111111111111111111111111111111111111111111111110110011111011010111111111001111111111111111111111111111111111111100111111111011010111111111111111110101111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111001111111111111111101100111111111111111111111111111111111111111111111111111111111101001111111100011111111111111111111111111111111111111111111111111110110011111110110011111111111111111111111111111111111111111111111111111011001111111111111111111111111110001111111111010111111111111111111111111111111111111111111111111111111111111111010111111010111111111111111111111111111111111011001111111010011111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111110111111110101111111111111111111111111111111111111011011111111111101101111111111111111111111111111111111111110011111111111011001111111011010111111111111111111111111111111110100011101100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000011111111110000000000000000000000000000000000000000000000001011111110000001111111111111111000000000000000001111000000000011111111111000000000101111111111111111111111111111111000000000001011111111111111111110000000000000000000000000000000000000000000011111111111111111111111111111111111111110000000000010111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111110110100111111101101001111111111111111111111111111111111111111111111111110110000111111101100111111111111111111111111111111111111111111111111111111101100111110110100111111110011111111111111111111111111111111111010101111111110110011111111111111111101001111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111110110011111111111111111011001111111111111111111111111111111111111111111111111111111110001111111111010111111111111111111111111111111111111111111111111111110101111110100011111111111111111111111111111111111111111111111111111111001111111111111111111111111111010111111111010111111111111111111111111111111111111111111111111111111111111111010111111011011111111111111111111111111111111101011111111101011111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111110011111110110111111010101111111111111111111111111111111111111010111111111111100011111111111111111111111111111111111110101111111111101100111111111101011111111111111111111111111111111011001110100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000111111110000000000000000000000000000000000000000000000001011111100000001111111111111111110000000000000000011000000000011111111110100000000011111111111111111111111111111111000000000001111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111101010111111110110011111111111111111111111111111111111111111111111111111010010111111011010111111111111111111111111111111111111111111111111111111010101111111101011111101100111111111111111111111111111111111111101011111111101101011111111111111111010111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111110101111111111111111111010111111111111111111111111111111111111111111111111111111110100111111111010011111111111111111111111111111111111111111111111111101100111111110101111111111111111111111111111111111111111111111111111111010111111111111111111111111110110111111111010111111111111111111111111111111111111111111111111111111111111111010111111010111111111111111111111111111111111010111111111101011111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111110101111111111011111111010111111111111111111111111111111111111101101111111111111010111111111111111111111111111111111111110101111111110110011111111101101111111111111111111111111111111111101011100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111000000000000000000000000000000000001010110000000000010111110000001111111111111111111100000000000000000000000000011111111111000000000011111111111111111111111111101000000000000101111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110110100111111101101001111111111111111111111111111111111111111111111111110110101111110110011111111111111111111111111111111111111111111111111111110101011111011010011111111001111111111111111111111111111111111111111111111111011001111111111111111110101111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111101011111111111111110110011111111111111111111111111111111111111111111111111111110110101111111100011111111111111111111111111111111111111111111111111101100111111101000111111111111111111111111111111111111111111111111111111001111111111111111111111111111010111111111010111111111111111111111111111111111111111111111111111111111111110110111111010111111111111111111111111111111111100111111111101011111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111011111111011011111111011111111111111111111111111111111111111101011111111111111001111111111111111111111111111111111111111111111111110110111111110110011111111111111111111111111111111101000110000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111000000000000000000000010010101010111111111100000000010111100000001111111111111111111111000000000000000000000000011111111111000000000101111111111111111111111110100000000000000011111111111111111111101000000001001010101010101010000000000000000000000011111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111101001111111110110101111111111111111111111111111111111111111111111111101101001111111101001111111111111111111111111111111111111111111111111111111111111111110100111111110011111111111111111111111111111111111111111111111110110011111111111111111101011111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111011001111111111111111110100111111111111111111111111111111111111111111111111111111101100111111101101111111111111111111111111111111111111111111111111111101011111101100111111111111111111111111111111111111111111111111111110110111111111111111111111111110110011111110110011111111111111111111111111111111111111111111111111111111111111010111111010111111111111111111111111111111111100111111111100111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111011011111111101011111111111111111111111111111111111111111111110110011111111111101011111111111111111111111111111111111111111111111111011001111111111001111111111111111111111111111111110100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000010111111111000000000000000011011111111111111111111111110000000010111110000000111111111111111111111110000000000000000000000011111111111000000000000111111111111111111111010000000000000001111111111111111111111110000000000111111111111111111101111000000000000000000011111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110110101111111101101011111111111111111111111111111111111111111111111111111010011111110110011111111111111111111111111111111111111111111111111111111111111111101001111111100111111111111111111111111111111111111111111111111101100111111111111111011010111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111010011111111111111111101011111111111111111111111111111111111111111111111111111101101011111101001011111111111111111111111111111111111111111111111111011001111111101011111111111111111111111111111111111111111111111111110110011111111111111111111111111110111111110100011111111111111111111111111111111111111111111111111111111111111010111111010111111111111111111111111111111101100111111101000111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111100111111111101111111111111111111111111111111111111111111111110101111111111101100111111111111111111111111111111111111111111111111111101011111111100101111111111111111111111111111101101000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000101101111111111100000000000000111111111111111111111111111111010000000010111100000000011111111111111111111111100000000000000000000011111111111000000000000111111111111111010000000000000000001011111111111111111111111110000000000111111111111111111111111101100000000000000000111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111101101001111111010110011111111111111111111111111111111111111111111111111110100111111101100111111111111111111111111111111111111111111111111111111111111111110100011111110101111111111111111111111111111111111111111111111111011001111111111111110110101111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111110101111111111111111011001111111111111111111111111111111111111111111111111111111101001111111101011111111111111111111111111111111111111111111111111111010111111010001111111111111111111111111111111111111111111111111111110011111111111111111111111111100011111110110011111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111101010111111101100111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111101010111111101101111111111111111111111111111111111111111111111010101111111111101101111111111111111111111111111111111111111111111111101101111111101100111111111111111111111111111111101000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001001111111111111111100000000000011111111111111111111111111111111010000000010111110000000011111111111111111111111111000000000000000000011111111110100000000000000011101110000000000000000000000011111111111111111111111111101000000001011111111111111111111111111111110000000000000001111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111110110101111111101100111111111111111111111111111111111111111111111111111010010111111111001111111111111111111111111111111111111111111111111111111111111111101000111110101111111111111111111111111111111111111111111111111110110011111111111111101101011111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111101100111111111111111111010111111111111111111111111111111111111111111111111111111111010111111110001111111111111111111111111111111111111111111111111111010111111011001111111111111111111111111111111111111111111111111111110101111111111111111111111111110101111110110101111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111101011111111101101111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111101101111111101011111111111111111111111111111111111111111111111110111111111110110111111111111111111111111111111111111111111111111110110011111111110101111111111111111111111111111111101000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001001111111111111111111110000000000001111111111111111111111111111111111010000000000101100000000011111111111111111111111111110000000000000000011111111111110000000000000000000000000000000000000000010111111111111111111111111111110000000000111111111111111111111111111111111110000000000000111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111101101001111111011010111111111111111111111111111111111111111111111111111110100111111110100111111111111111111111111111111111111111111111111111111111111111010001111111111111111111111111111111111111111111111111111111111101010111111111111111011001111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111101011111111111111111110101111111111111111111111111111111111111111111111111111111010011111111010111111111111111111111111111111111111111111111111110110011111111010111111111111111111111111111111111111111111111111111101101111111111111111111111111110101111111110101111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111101101111111110101111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111110011111110101111111111111111111111111111111111111111111111101011111111111111010111111111111111111111111111111111111111111111111111010111111111010111111111111111111111111111111110110010100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111110000000000001111111111111111111111111111111111010000000000101110000000011111111111111111111111111111100000000000000011111111111110000000000000000000000000000000000000001011111111111111111111111111111110000000000111111111111111111111111111111111111110000000000011111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110110011111111110100111111111111111111111111111111111111111111111111111101001111111011011111111111111111111111111111111111111111111111111111111111111110100101111111111111111111111111111111111111111111111111111111111011011111111111111110110011111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111010111111111111111101101111111111111111111111111111111111111111111111111111111100011111111100011111111111111111111111111111111111111111111111111110011111110100011111111111111111111111111111111111111111111111111101101111111111111111111111111110101111111110101111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111101011111111110101111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111110110111111110101111111111111111111111111111111111111111111111111011111111111011001111111111111111111111111111111111111111111111111011011111111010101111111111111111111111111111111111001111110000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111010000000000101100000000111111111111111111111111111111110000000000000011111111111111100000000000000000000000000000000000101111111111111111111111111111111110000000000111111111111111111111111111111111111111110000000011111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111101101001111111011010111111111111111111111111111111111111111111111111111010101111110101111111111111111111111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111111111111110110111111111111111101000111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111110110011111111111111111101011111111111111111111111111111111111111111111111111111101000111111110101111111111111111111111111111111111111111111111111101101111111110011111111111111111111111111111111111111111111111111101101111111111111111111111111101001111111110101111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111101011111111110011111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111001111111110101111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111101100111111101100111111111111111111111111111111111010111111111100000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000101111111111111111111111111111111111110100000000101110000000111111111111111111111111111111111110000000000011111111111111111000000000000000000000000000001011111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111001111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111",
"0111111111111111111111111111111111111111111111111111111111111111111111111111111010011111110110100111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111101100111111111111111011001111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111101100111111111111111011001111111111111111111111111111111111111111111111111111101101011111101100111111111111111111111111111111111111111111111111101100111111110100111111111111111111111111111111111111111111111111111100111111111111111111111111101100111111110101111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111101011111111110011111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111001111111011011111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111110101111111110101111111111111111111111111111111101010111111101100000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000010111111111111111111111111111111111111110100000000011111100011111111111111111111111111111111111111110000111111111111111111111110000000000000000000000010111111111111111111111111111111111111111101000000101111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111",
"0010011111111111111111111111111111111111111111111111111111111111111111111111111101101011111111010001111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111011011111111111111111010011111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111101011111111111111110110111111111111111111111111111111111111111111111111111111010011111111101011111111111111111111111111111111111111111111111111101011111101101111111111111111111111111111111111111111111111111111010111111111111111111111111101000111111101101111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111101011111110110011111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111011011111111101111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111010111111110110011111111111111111111111111111110101011111111110001010000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100001111111111111111111111111111111111111111111111111111111111111111111111111111111111010000010001010111111111111111111111111111111111111111111111101000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1000001011111111111111111111111111111111111111111111111111111111111111111111111111011010011111110110100111111111111111111111111111111111111111111111111110001011111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111110101011111111111111110100111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111011001111111111111111110011111111111111111111111111111111111111111111111111111011010111111110001111111111111111111111111111111111111111111111111011011111111000111111111111111111111111111111111111111111111111111010111111111111111111111111111100111111101100111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111101111111110110011111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111100111111101011111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111011111111111001111111111111111111111111111111110101111111110100000111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101100010011111111111111111111111111111111111111111111111111111111111111111111111111101100111111111011001111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111101011111111111111111101001111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111110110011111111111111101100111111111111111111111111111111111111111111111111111110100111111111010111111111111111111111111111111111111111111111111111001111111101011111111111111111111111111111111111111111111111111011011111111111111111111111111101011111101100111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111100111111110011111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111101011111111011011111111111111111111111111111111010111111111010000011101000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111110100001001111111111111111111111111111111111111111111111111111111111111111111111111111010011111110110010111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111010101111111111111111010111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111110101111111111111111101011111111111111111111111111111111111111111111111111111110101111111110011111111111111111111111111111111111111111111111110101111111011001111111111111111111111111111111111111111111111111111011111111111111111111111111101011111101100111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111101011111110110111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111101101111111101101111111111111111111111111111111111011111111111100001110100001001000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111011000011111111111111111111111111111111111111111111111111111111111111111111111111110100111111101101011111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111111111111111111111111111111111110101111111111111111110101111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111101100111111111111111111001111111111111111111111111111111111111111111111111111101001111111110101111111111111111111111111111111111111111111111110110111111111001111111111111111111111111111111111111111111111111111001111111111111111111111111011011111111101011111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111110011111110101111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111110011111110110011111111111111111111111111111111101111111111110000111111000101111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110110001001111111111111111111111111111111111111111111111111111111111111111111111111011010011111110110010111111111111111111111111111111111111111111111110100011111111111111111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111010011111111111111110110011111111111111111111111111111111111111111111111111111101011111101100111111111111111111111111111111111111111111111111110011111111010111111111111111111111111111111111111111111111111110101111111111111111111111111010011111111101011111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111110110111111111011111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111010111111111010111111111111111111111111111111110111111111110100011111100000111111010000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1001111111111111011000011111111111111111111111111111111111111111111111111111111111111111111111110101100111111101100101111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111010111111111111111110101111111111111111111111111111111111111111111111111111010011111111101011111111111111111111111111111111111111111111111101011111111100011111111111111111111111111111111111111111111111110101111111111111111111111111011011111111101011111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111110110111111010111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111011011111111011011111111111111111111111111111111011101111111010010111101001011111111110100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010100111111111110101001001111111111111111111111111111111111111111111111111111111111111111111111111011010111111111010111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111010010111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111110011111111111111101100111111111111111111111111111111111111111111111111111111010111111011001111111111111111111111111111111111111111111111101010111111110011111111111111111111111111111111111111111111111110110111111111111111111111111011001111111101011111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111011001111111010111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111101100111111101100111111111111111111111111111111101011111111101101011110100100111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101101001111111111111111000101111111111111111111111111111111111111111111111111111111111111111111111111110100111111101100101111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111101001111111111111111011001111111111111111111111111111111111111111111111111110100111111111010111111111111111111111111111111111111111111111111010111111110101111111111111111111111111111111111111111111111111101011111111111111111111111111001111111010111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111011011111101101111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111110101111111110011111111111111111111111111111111101111111111110100111111010011111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111010101111111111110101101001111111111111111111111111111111111111111111111111111111111111111111111111011001111111111010011111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111011011111111111111111010111111111111111111111111111111111111111111111111110110101111110100011111111111111111111111111111111111111111111111010111111101100111111111111111111111111111111111111111111111110101011111111111111111111111111010111111011011111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111010111111101011111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111010111111110101111111111111111111111111111111110111111111110110011111101011111111111111111111000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111101001111111111111011010101111111111111111111111111111111111111111111111111111111111111111111111110110100111111101100111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111011001111111111111110110011111111111111111111111111111111111111111111111111101100111110110011111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111101011111111111111111111111111010111111011001111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111101010111111101011111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111001111111011001111111111111111111111111111111011111111111011001111110100111111111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110110100111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111011001111111011010111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111110100011111111111111101101111111111111111111111111111111111111111111111111111101011111101101111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111101011111111111111111111111110110111111111011111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111101011111111101111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111101011111111010111111111111111111111111111111111011111111101101011110110101111111111111111111111010000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111011001111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111110110100111111101100111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111101101111111111111111101011111111111111111111111111111111111111111111111111010001111111100111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111101011111111111111111111111110110011111111001111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111110111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111101101111111101011111111111111111111111111111111101111111111110101111011010111111111111111111111111011000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111110101011111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111101010111111011001111111111111111111111111111111111111111111111101001011111111111111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111100111111111111111011011111111111111111111111111111111111111111111111111111010111111011011111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111011111111111111111111111110110011111110101111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111110111111111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111110110011111111101011111111111111111111111111111110111111111111010011101101011111111111111111111111111110000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111011001011111111111110110011111111111111111111111111111111111111111111111111111111111111111111111110110101111110101101111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111011001111111111111111001011111111111111111111111111111111111111111111111110100011111011001111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111110110011111110101111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111010111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111001111111110111111111111111111111111111111111111111111111010101110110101111111111111111111111111111011000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1011111111111111111111111110100111111111111111011001111111111111111111111111111111111111111111111111111111111111111111111101101001111111011001111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111010001111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111010111111111111111110011111111111111111111111111111111111111111111111111110101111110110111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111111110101111110111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101111111011111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111011001111111010111111111111111111111111111111111011111111101011111111010111111111111111111111111111111010000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010100111111111111111111111111010011111111111110110100111111111111111111111111111111111111111111111111111111111111111111111110110101111110101010111111111111111111111111111111111111111111111011001011111111111111111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111110011111111111111101101111111111111111111111111111111111111111111111111101100111110110011111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111101100111111101011111111111111111111111111111111111111111110110111111011001111111111111111111111111111101000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101101010111111111111111111111101100101111111111111011001111111111111111111111111111111111111111111111111111111111111111111111101101001111111010111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111101100111111111111111100111111111111111111111111111111111111111111111111111100111111101101111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110101111111111111111111111111111111111111111111111001111101100111111111111111111111111111110100000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111110110100111111111111111111111110110011111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111010101111110101111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111101001111111111111111001111111111111111111111111111111111111111111111111011001111101100111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111110101111111111111111111111111111111111111111111100101110110011111111111111111111111111111010010100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111101101010111111111111111111111101101001111111111111011001011111111111111111111111111111111111111111111111111111111111111111111101101001111111011111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111010111111111111110101111111111111111111111111111111111111111111111111111001111111010111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111011111111111111111111111111111111111111111111101101111110101111111111111111111111111111101001001010000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110110010101111111111111111111110110101111111111111110100101111111111111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111110110011111111111111110011111111111111111111111111111111111111111111111110110111111011001111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111110110011111100111111111111111111111111111110100100111010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010101010101010101001011111111111111111111111111111111111111111111111111111111010101010101001011111111111111111111111111111111111111111111111111111111110100000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111011010010111111111111111111111011001011111111111010101011111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111110100111111111111101101111111111111111111111111111111111111111111111111110101111110101111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111101101111111101011111111111111111111111111111111111111111011001111101101111111111111111111111111111110010011111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010000000000000000000000000001010101111111111111111111111111111111111111111111010100000000000000000001010111111111111111111111111111111111111111111111111101000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111101101011111111111111111111110101100111111111111101100111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111101011111111111111011011111111111111111111111111111111111111111111111101100111110101011111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111101100111110110011111111111111111111111111101100001111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101000000000000000000000000000000000000000000011111111111111111111111111111111111110100000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111010110011111111111111111111111011010111111111111010110011111111111111111111111111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111011001111111111111010101111111111111111111111111111111111111111111111111101011111101011111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111110101111011011111111111111111111111111111110000111111110000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000111111111111111111111111111111101000000000000000000000000000000000000010111111111111111111111111111111111111101000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111101101001111111111111111111110101100111111111111101101011111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111010111111111111110101111111111111111111111111111111111111111111111111011001111111011111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111110110111101100111111111111111111111111111110110011111110100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000000000000000000000000001111111111111111111111111101000000000000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000000000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111110110100111111111111111111111010101011111111111010110011111111111111111111111111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111111111101011001111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111110101111111111111101011111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111011001111101011111111111111111111111111111100001111111011000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000101011000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111011010111111111111111111111101010111111111111101101011111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111101100111111111111111011111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111101100111110110111111111111111111111111111101101011111101100000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001001010101010101010101010101010000000011111111111111111101000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000001011111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111101100111111111111111111111110101011111111111110110011111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111111111111111111111101010111111111111111111111111111111111111111111111010011111111111111010111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111110101111011011111111111111111111111111110100101111011000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000001001011111111111111111111111111111110100000000111111111111110100000000000000000000010101010101010101100000000000000011111111111111111111111110000000000000000111111111110100000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111011001011111111111111111111101010101111111111111101001111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111111111111111111111101011011111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111001111111100111111111111111111111111111010001111101000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111100000000111111111111111000000000000000010101111111111111111111110101000000000000111111111111111111111000000000000000011111111111111000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111101100101111111111111111111110110011111111111110110010111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111011011110101011111111111111111111111111101101011111101000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000111111111111111111111111111111111111100000000111111111111010000000000000101111111111111111111111111111111110000000000111111111111111111100000000000000001111111111111110100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111010011111111111111111111111011001111111111101101001111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111101100111111001111111111111111111111111110110100111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111100000000111111111101000000000010111111111111111111111111111111111111111000000000011111111111111111100000000000000111111111111111111101100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111011001111111111111111111110110101111111111110110100111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111110110011111100111111111111111111111111111111010011111111111100000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111110000000000111111110100000000001011111111111111111111111111111111111111111100000000001111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110101010111111111111111111111011001111111111111010101111111111111111111111111111111111111111111111111111111111111111111010001011111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111001111101011111111111111111111111111111101001111111111110101000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111110000000000111111111000000000101111111111111111111111111111111111111111111100000000001111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111010101111111111111111111111101100111111111110101100111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111110101100111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111100111111010011111111111111111111111111110100111111111110101110100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111111111111111000000000000111111010000000010111111111111111111111111111111111111111111111100000000001111111111100000000000000111111111111111111111111111111111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111101100111111111111111111111011010011111111111010110111111111111111111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111101101111010101111111111111111111111111111010011111111111101011111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111111111111100000000000000111101000000001011111111111111111111111111111111111111111111111100000000001111111111100000000000011111111111111111111111111111010101010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111101100111111111110101010111111111111111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111110110011111011111111111111111111111111111100111111111111110001111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111111111111100000000000011111111000000001111111111111111111111111111111111111111111111111100000000001111111101000000000000011111111111111111110101010110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111101100101111111111111111111010110011111111111010101011111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111011001111110011111111111111111111111111101100111111111111000011111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111111111010000000000000011111110000000011111111111111111111111111111111111111111111111111100000000001111111110000000000001111111111111010101100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111001010111111111111111111101101001111111110101010111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111100111111010111111111111111111111111110110011111111111100001111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111111111100000000000001111110100000000111111111111111111111111111111111111111111111111110100000000001111110100000000001011111111111110000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111101011001111111111111111111110110011111111111011010011111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111110101111011011111111111111111111111111011001111111111110000111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111111101100000000000001111111100000010111111111111111111111111111111111111111111111111110000000000001111111000000000000111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111111111101011001111111111101010111111111111111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111110110111111100111111111111111111111111101010111111111111000011111111111111111111000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111100000000000000111111111000000000111111111111111111111111111111111111111111111111110000000000101111010000000000101111111111111100000000000000000000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111110110100111111111110101111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111010101011111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111011001111110111111111111111111111111111110011111111111100010111111011111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111010000000000000011111111110000000001111111111111111111111111111111111111111111111111010000000000111111010000000000011111111111111110000000000000000000000000000010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010101111111111111111111011001111111111101011111111111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111100111111001111111111111111111111111111001111111111110101011111111111111111111110100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111000000000000001001111111110000000011111111111111111111111111111111111111111111111111000000000000111111010000000010111111111111111111100000000010101001000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111110100111111111111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111110101111011011111111111111111111111111100101111111111000101111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111110100000000000000101111111111110000000010111111111111111111111111111111111111111111111101000000000010111101100000000010111111111111111111111001100111111101000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111010110011111111111111111111111111111111111111111111111111111111111111111111111111111010110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111110110111101011111111111111111111111111101011111111111010001111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111110000000000000010011111111111110000000000111111111111111111111111111111111111111111110100000000000011111111000000000001111111111111111111111111111111111110000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111011011111111011111111111111111111111110110111111111110000111111111111111111111111111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111000000000000001011111111111111110000000010111111111111111111111111111111111111111111111000000000001011111101000000001011111111111111111111111111111111110100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111101100111111111111111111111111111111111010101111111110110011111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111100000000000000001011111111111111110000000000101111111111111111111111111111111111111111010000000000001111111111000000000011111111111111111111111111111111010000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111111111101101011111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111101011111111111111111111111111111111101011111111111011001111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111110000000000000000101111111111111111010000000000101111111111111111111111111111111111111110000000000000011111111101000000001011111111111111111111111111111101000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111110101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111001111111111111111111111111111111110101111111111101000111111111111111111111111111111111111111100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111100000000000000000010111111111111111111110100000000001011111111111111111111111111111111010000000000000010111111111111000000001011111111111111111111111111111101000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111010101111111111111111111111111111111110111111111110110101111111111111111111111111111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000101111110000000000000000001001111111111111111111111100000000000000101111111111111111111111110100000000000000000001111111111101000000001011111111111111111111111111010000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111011000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000100111111111111111111111110100000000000000001011111101111111110100000000000000000000000111111111111111000000000011111111111111111111111101000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011001111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111010000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111101000000000000000000000000000000000000000000000000000000011111111111111101000000000010111111111111111111110100000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101010111111111111111010110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111010000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001011111111111111111111111111111111010000000000000000000000000000000000000000000000000010111111111111111111000000000010011111111101110100000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101011010011111111111111101101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111011001011111111111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111100101111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111011000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000100111111111111111111111111111111111010000000000000000000000000000000000000000000000000111111111111111111101000000000000001001010100000000000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111101101001111111111111110101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111110000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000010111111111111111111111111010000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110110100111111111111111010110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101011111111111111111011001011111111111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111110101101111111111111111111111111111111111111111111111111111111000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000101111111111111111111111111111111111111111111101000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111011010010111111111111101011001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101111111111111111101100101111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000001011111111111111111111111111111111111111111111111111011000000000000000000000000000000010111111111111111111111111111111111100000000000000000000000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111110101101001011111111111110110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101011111111111111111111010011111111111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111101010111111111111111111111111111111111111111111111111111111111111000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000010111111111111111111111111111111111111111111111111111111111101100000000000000000000010101111111111111111111111111111111111111101000000000000000000000000001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111110110100111111111111111110101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111101101010101010101111111111111111111111111111111111111111111111111000000000000000001010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111101010101011111111111111101011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111110100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101101001011111111111110101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111101001011111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111110101100111111111111111110110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111110100001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111011010010111111111111101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111011001011111111111111111111111111111111111111111111111111111111111111111111101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111101011001011111111111111101011001111111111111111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111110110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111110110010101111111111111010110100111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111110101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110101010111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111101000111111111111111111111111111111111111111111101100000000010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111110100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111101010101111111111111111101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111010011111111111111111111111111111111111111111111111111111111111111111111101011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111110001011111111111111111111111111111111111111110110001010101000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111110110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110101011101111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111011001011111111111111111101001111111111111111111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111110001011111111111111111111111111111111111111110100000111111111011000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111101111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111101010010111111111111111111111111110010111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111101101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010111110000000000001011111111111111111111111111111111111111101000111111111111111111111111111111111111111111111111111111111111111111111111101011001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111101011011111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110100000101101000000111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111101101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111110110010101111111111111010110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100000011111110110000010011111111111111111111111111111111000101111111111111111111111111111111111111111111111111111111111111101011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111011001010111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111110100000010111111111111011000001001111111111111111111111111011000111111111111111111111111111111111111111111111111111111111111011001011111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111100001111111111110000001111111111111111101000010111111111111111111111111100001111111111111111111111111111111111111111111111111111101011001100101111111111111111111010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111101000010111111111110000011111111111111111111011010111111111111111111111101001001111111111111111111111111111111111111111111111111010110010111111111111111111101010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111100010011111110100000001111111111111111111111111111111111111111111111101000111111111111111111111111111111111111111111111010110100101111111111111111111010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111010101010101010101011101111111111101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111000000101100010010000111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111010110011001111111111111111101010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010110101010000000100000000000000000001010101010101010101010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111110110000000001011111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101001111111111111111111010110010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010101000000000000000000000000000000000000000000000000000000000000000000010001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100011111111111111111111111111111111111111111010101011111111000101111111111111111111111111111111111111111111111111111111111111111111111111111110101101001011111111111111101010110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010110101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010101010100111111111111111111111111111111111111111111111101010101010101010011111111111111111111111111111111111110110101010100000000000111111111111111111111111111111111111111111111111111111111010101010101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111100101111111111111111111111111111111111111111111111111111111111111111111111111101011001011111111111111101010110010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010011111111111111111111111111111111111111111111111111000000010111111111111111111111111111111111111111101101010101010001011111111111111111111111111111111111111111111111010101010000000000000000111111111111111111111111111111111111111101010000000000000000000000111111111111111111111111111011010100000000000000000000000101111111111111111111111111111111111111111111111110110100000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011001011111111111111101011010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101000000000000000000000000000000000000000100000000010100110001001010101000000000000000000000000000000000000000000000010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111000100010111111111111111111111111111111110000000000111111111111111111111111111111111111100000000000000000000000001011111111111111111111111111101000100010000000000000000000000000000111111111111111111111111111111111111010000000000000000000000000001011111111111111111111111000000000000000000000000000000000101111111111111111111111111111111111111111111101100000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111110101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111101011010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000000000000000000000001010010101010111010110100111111110001011111111000001011010000000000000000000000000000000000000000000101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000011111100000000000111111111111111111111111111111110000000000101111111111111111111111111111110000000000000000000000000000000000111111111111111111010010000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111111111011000000000000000000000000000000001111111111111111111111111111111111111110110000111111111111111111111111111111111111111111111",
"1111111111010101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111101011001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100000000000000000000000000000000000101010011111111111111111111111111111010111111111101011111111100001110101000000100000000000000000000000000000001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000011111000000000000001111111111111111111111111111110000000000001111111111111111111111111110000000000000000000000000000000000000001011111111111110000000000000000000000000000000000000000000000111111111111111111111111111010000000000000000000000000000000000101111111111111111110000000000000000000000000000000000100101111111111111111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111111100000000000010111111111111111111111111111111111111111111",
"0111111111111111011010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000000000000010001000100010001000000000000010110110101111111101101111111111011111111111111111011111111111011001010110000000000000000000000000000000001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010011111000000000000001111111111111111111111111111110000000000011111111111111111111111110000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000101111111111111111111111110100000000000000000000000000000000000000111111111111111111000000000000000000000000000010010101111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111111111000000000000000010111111111111111111111111111111111111111111",
"0010011111111111111111010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010000000000000000000000000011111110111111101111101010101101000011110101111111110000111111101000111111111100111111111011111111111111101011010000000000000000000000000000000001010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000111111000000000000001111111111111111111111111111110000000000111111111111111111111111000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000001001111111111111111111111111010000000000000000000000000000000000000011111111111111111111000000000000000000000000100111111111111111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111000000000000000000000010111111111111111111111111111111111111111111",
"1000001010011111111111111101011001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101000000000000000000000000010100001111111010010111111110110111111110101011111111111111101111111111101100111111101001011111111100001111111011001111101010000000000000000000000000000000000001010101010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111000000000000000011111111111111111111111111110000000000111111111111111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001110111011111111111111111111111111101000000000000000000000000011101110110001111111111111111111111000000000000000000100111111111111111111111111111111111111111111111111111110000000000000000000000001011011101110001111111111111111111111111110000000000000000000000000010111111111111111111111111111111111111111111",
"0110100000001010011111111111111101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010000000000000000000000000100010111111010101111111111010111111111000011111110100011111111110011111111101011111111111111101100101111101101011111111010001111111010000010101100000000000000000000000000000000000000000100010101001010111010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000101111000000000000000011111111111111111111111111110000000000111111111111111111000000000000000000000011111111011111011100000000000000001111111111100000000000011100000000000011111111111111111111111111111111010000000000000000000000011111111111111111111111111111111111111111000000000000001011111111111111111111111111111111111111111111111111111100000000000000000000001011011111111111111111111111111111111111111000000000000000000000000000100111111111111111111111111111111111111111111111",
"1111010110100000001001111111111111111101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000010100111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101101000000000000000000000000000000010011111101011111111110111111111111111110101111111110110011111110100101111111110000101010110101000000000000010000111111111110111111111111001111111011000010110100000000000000000001010100000000000000000000000100000100010101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111000000000000000000111111111111111111111111110000000000111111111111111111000000000000000011111111111111111111111111110100000000000011111111111111111101111100000000001011111111111111111111111111111111010000000000000000101111111111111111111111111111111111111111111111110000000000100111111111111111111111111111111111111111111111111111111100000000000000001011111111111111111111111111111111111111111111100000000000000000000000001011111111111111111111111111111111111111111111111111",
"1111111111110110100000100111111111111101110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101000000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000000000000000000000000000000000010101011111111101001111111101001111111111001111111110101111111111111111101011101011000000000000000000010101010000000001011101001111111110111111111111111111111111111011010100110100000011111110110000101011000000000000000000000000000000010101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000101111000000000000000000111111111111111111111111110000000000111111111111111100000000000000111111111111111111111111111111111111000000000011111111111111111111111100000000001111111111111111111111111111111101000000000000000001111111111111111111111111111111111111111111111111010000000000111111111111111111111111110111011101111111111111111111110000000000000000100111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111",
"1111111111111111110110000000010111111111111111011101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010100000101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011000000000000000000000000000000010100000000111111111111111010111111111011001111111010010111111111000111111110110010101101000000010101001100111011111111111100111011111101011111111100001111111111010111111110101111111111111010101111111111101010111111101000101011000000000000000000000000000000010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101100000000000000000000001111111111111111111111110000000000111111111111110000000000001111111111111111111111111111111111111111000000001001111111111111111111111100000000001111111111111111111111111111110100000000000000101111111111111111111111111111111111111111111111111111000000000000111111111111111111010101000000000000111111111111111111000000000000000011111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111110110000010101111111111111111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010100000000000000000000000000000101000100111110110000111111111100111111111010111111111110111110111111111111001011111011000000000101000100111111110101111111101011111111111111111110111111111011011111111010010111111111000011111110100011111111101011111111111011111111111111111101000000000000000001000000000000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000101100000000000000000000000111111111111111111111110000000000111111111111100000000000111111111111111111111111111111111111111111110000000010111111111111111111111100000000001111111111111111111111111111010000000000000010111111111111111111111111111111111111111111111111111111000000000000111111111111011101000000000000000010111111111111110100000000000000001111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111011000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101000000000000000000000000000000000100101111101011111111101100111111101001011111111100011111111011011111111110101111111010110100010100111110110011111110110101111111101000111111101101011111111010111111111110111111111111111111001111111111010011111110100101111111110101111111101010111111101100000000000100101011010000000000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101110000000000000000000001011111111111111111111110000000000111111111111000000000011111111111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111111000000000000001011111111111111111111111111111111111111111111111111111111000000000010111111110101000000000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101011010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010110000000000000000000000000101010000000001001110110011111111101011111111111111111011111111111100111111111100001111111010010010110000000100101110101111111111111111101111111111101101111111101101011111111100011111111011001111111110101111111111101111111111111111101011111111110100111111110000111111101000001100000001001111111011010000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101110000000000000000000000001111111111111111111110000000000111111110100000000001111111111111111111111111111111111111111111111010000000010111111111111111111111100000000001111111111111111111111111101000000000000101111111111111111111111111111111111111111111111111111111111000000000000111101010000000000000000000000000011111111111111011000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111101101000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101010000000000000000000100001010111010110001010111111110110101111111110101111111101100111111111011111111111011111110111111111010000101010011010111111111000011111110110101111111101011111111111011111111111111111010111111111100001111111010010111111111010111111110110111111111101111111111111111111010111111111100111110110000000010111011001011010000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111000000000000000000000010111111111111111111110000000000111111111000000000111111111111111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111100000000000010111111111111111111111111111111111111111111111111111111111111000000000000101000000000000000000000000000001011111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111110101100010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110100000000000000000000010010111011001111101100000100111111111111101111111111110101111111110000111111101000111111111101011111111010101100010010111110101111111110110111111110110011111111100100111111110100111111101010111111111011111111111111111110101111111111010111111111000011111110110101111111101101111111111011111111111111111010000001001010001111111010000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111000000000000000000000000011111111111111111110000000000111111111000000001111111111111111111111111111111111111111111111111110000000010111111111111111111111100000000001111111111111111111111111100000000000011111110100110101001101010011010100101111111111111111111111111000000000000000000000000000000000000001010111111111111111111100000000000111111101001101010011010100110100110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111110110100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010001000000000000000101001101001111111100010011000000010111111111010011111111101011111111111111111011111111101100111111101101011111101100010100111011010111111110101111111111101111101111111111101011111111101000111111101001011111111101011111111011011111111110111110111111111111101111111110110101111111110100111111110000111111101100111111110000000101111111111110101100000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000100111000000000000000000000000101111111111111111110000000000111111011000000011111111111111111111111111111111111111111111111111110000000000111111111111111111111100000000001111111111111111111111111100000000000010100000000000000000000000000000000000101001111111111111111111000000000000000000000000000000001010101111111111111111111111000000000000101010000000000000000000000000000000001010011111111111111111111111111111111111111010101010101010101010101010101010101010101010101001111111",
"1111111111111111111111111111111111111111111111111111110110100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000100110101111111111111111111010000010011001111111111010011111111000011111111110101111111101011111111111111111011111010110001001111111010001111111110010111111111010011111111110011111111111111111111111111101010111111111101011111111100001111111010001111111111001111111110111111111111111111101011111111101101111111101001011111111000000000101011001111111011000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111000000001000000000000000000111111111111111110000000000111111100000000111111111111111111111111111111111111111111111111111100000000010111111111111111111111100000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000100111111111111111000000000000000000000000000000101111111111111111111111111111010000000000000000000000000000000000000000000000000000001010111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111",
"1111111111111111111111111111111111111111111111111111111111010110001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000000000000000000001011111101001011111111101001011000000011111111111111111101111111110110011111111110101111111110000111111101000111111101100010111111111111111111111111110101111111111010011111110100011111111100101111111101101111111111011111111111111111010111111111011001111111111010111111111000011111110110011111111101011111111111111111010111111111011010000010000001111111010010011000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111000000001110000000000000000001111111111111110000000000111111010000001011111111111111111111111111111111111111111111111111000000000000111111111111111111111100000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000100111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000101111111111111111111111111111100000000000000000000000000000000000000000000000000000101111",
"1111111111111111111111111111111111111111111111111111111111111111011000001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000000000100101111111111111100111111111100000001010100001111111011010111111110101111111111111111101111111111101101111111101000111010000000011111111101001111111010101111111110111111101111111110101011111110110101111111110100111111101000111111111100111111111011111111101111111110101111111110110011111110100101111111110101111111101100111111111010111111111100000000011111111111001111111101000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111101000000101111000000101111000000000000000010111111111111110000000000111101000000001011111111111111111111111111111111111111111111111111000000000001111111111111111111111100000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000001011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000011111",
"1111111111111111111111111111111111111111111111111111111111111111111111011010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101000000000000010101000001111111101011111111111111111100000011111010101111111011010111111111000011111110100011111111101011111111111111111110110001001010111111111011001111111010001111111011010111111110110111111111101111111111111111101011111111101100111111101101011111111100011111111011001111111110101110111111111111101111111111110101111111110001111111101000111111111100000000010010101111111111111110101000000000010100111111111111111111111111111111111111111111111111111111111111111111111111101100000011111000000111111100000000000000000011111111111110000000000111101000000101111111111111111111111111111111111111111111111111100000000000011111111111111111111111100000000001111111111111111111111111111010000000000000000000000000000000000000000000000000000000000011111111111000000000000000001111111111111111111111111111111111111111111110100000000000000000000000000000000000000000000000000000000001011111111111111111111111111111010000000000000000000000000000000000000000000000000011111",
"1111111111111111111111111111111111111111111111111111111111111111111111111101101000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101000000000000000100111111110101111111110000111111101101010001011010111111111111111110111111111110101111111110110011111110100101111111110001111100000000111111111111111110111111111111011111111111010111111111010011111110100011111111110011111111101111111111111111111010111111111011001111111010001111111011010111111111010111111111101011111111111111101111111111101100111111111001001100000001001111111011001111111011000000000000010011111111111111111111111111111111111111111111111111111111111111111111101000000011111000000011111111000000000000000000111111111110000000000111110000000101111111111111111111111111111111111111111111111111100000000000011111111111111111111111100000000001111111111111111111111111111111000000000000000000000000010010100000000000000000000000000011111111111000000000000001111111111111111111111111111111111111111111111111101000000000000000000000000000101000000000000000000000000000011111111111111111111111111111111010101010101010101010101010101010101010101010111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111101101000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000000100111111111111101111111111101011111111101000000011111000011111111010001111111110101111111111101111101111111111101011111111110001000100110001011111101001011111111011011111111110111111111111111110101111111110110011111111100101111111110001111111101100111111111010111111111111111110111111111111010111111111000100111110100011111111110101111111101011111111111111111110111110100000001111111010010111111110000011000000000001001111111111111111111111111111111111111111111111111111111111111111101000000011111000000111111111110000000000000000001111111110000000000111101000000000111111111111111111111111111111111111111111111110000000000001111111111111111111111111100000000001111111111111111111111111111111101100000000101010101010111111101010101010110000000000000101111111111000000000001111111111111111111111111111111111111111111111111111111010100000001010101010101111111110101010101010000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000000000010100000011111110110011111111110011111111111110110001011111111010111111111011001111111010010111111111010011111110110111111111111111101100010111101001011111111100111111111100011111111010001111111011001111111110101111111111111111101111111111101101111111101000111111101101011111111101011111111110111111111111111110110001011110110011111110110101111111110000111111101100101111111010101100000011111111111111111110101110101100000000000100101111111111111111111111111111111111111111111111111111111111110000000111111000000011111111101000000000000000001111111110000000000111110000000000111111111111111111111111111111111111111111111000000000000001111111111111111111111111100000000011111111111111111111111111111111111110101111111111111111111111111111111111111011000000000011111111111000000000011111111111111111111111111111111110100000010111111111111111101010111111111111111111111111111111111110101000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000010100101110101111111110100011111111100101111111110001000011111100111111111111111110111111111110111111111111010111111110100011111110100101110100110101110101111011111111111111111010111111111011001111111110010111111111010011111110110011111111101111101111111111111011111111111100111111111100001111111010001111111011010111101000001111111111111111111111111111101101111111101000111111101001011111000001001111111111011111111111111010110000000000010011111111111111111111111111111111111111111111111111111111101000010111111000000111111111111010000000000000000011111110000000000111101000000001011111111111111111111111111111111111111111111000000000000111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111000000000011111111111111111111111111111100000000000010111111111111111111111111111111111111111111111111111111111111000000001011111111110000000001111111111111111111111111111111111111111111111111111111111111111111",
"0110101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111101000010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101110111111111111111111111111111111111111111111101000000000000000101110101111111111101111111111111111101011111110110001011111101000111111101101011111111011011111111110111111111111111110101111111110110011111011110001010011110000111111111100111111111011111111111111111111111111111111010111111110100011111110100101111111101100111111111011111111111111111011111111111011001111111011010111111010000011111110110011111110101011111111111111111111111111111010111111101000001111111010010111111011010111111011000000000001001111111111111111111111111111111111111111111111111111110000010111111000000011111111111111000000000000000000111110000000000111110000000000001111111111111111111111111111111111111111100000000000000111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000011111111111000000000011111111111111111111111100000000000000000010111111111111111111111111111111111111111111111111111111111100000000001011111111100000000000111111111111111111111111111111111111111111111111111111111111111111",
"1111110110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111011000001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111010101101010101010100010101000001000100010101001010111111111111111111111110110101000000000000001011111110010111111111010011111110101011111111111011000010111111101010111111111101001111111100001111111011010111111110101111111111101111111111111111101000001111101101111111101001011111111101011111111011001111111110111111111111111111111111111111110011111111110101111111110000111111111101011111111010111111111111111111111111111111000011111110100011111110100101111111110100111111111010111111111111111010000011111010111111111111010111111111000000000000010011111111111111111111111111111111111111111111111111110000010111111000000111111111111111110000000000000000001110000000000111101000000000010111111111111111111111111111111111111110000000000000011111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111101000000000010111111111111000000000011111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000001111111111100000000000000111111111111111111111111111111111111111111111111111111111111111",
"1111111111110110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110010111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111110000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101010100010001000000000000000000000000000000000000000000000000000000000000000100101111111011101101000000000000010011111111111111001111111111010011111110100101111111100001011111101101111111111111111111111111111110111111111011010111111110010011111111000011111110110011101101001011111111111111111111111111111011011111111100001111111010010111111111010111101111101111111111111111101011111111101010111111101001011111111100011111111011001111111110101110100000111111111111111111101011111111110100111111110000111111101101011110110001011111111110111111111111111110101010100000000001001111111111111111111111111111111111111111111110100000001111111000000011111111111111111100000000000000000010000000000111111100000000000010111111111111111111111111111111100000000000000001111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111110100000000000001111111111111000000000011111111111111000000000000000000000000001011111111111111111111111111111111111111111111111111111101000000000000101111111111110000000000000001111111111111111111111111111111111111111111111111111111111111",
"1111111111111111010110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101011111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101011000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010100000000000000000001001111111011011111111111111111111111111110101111111011000011111111110001111111101000111111111100111111111010111111111111111110101111111110110111111110100101110101110101111111101100111111111010111111111111111111111111111011001111111111010111111111000011111110110101111111101011111111111111111111111111111100111111111100001111111010010111101000010011111110101011111111111011111111111111111011111111101100111111111000010111111010001111111011001111111111110100000000000011111111111111111111111111111111111111111110110000001111111000000111111111111111111111000000000000000000000000000111111100000000000000001111111111111111111111101100000000000000000001111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111110101000000000000000111111111111101000000001111111101110000000000000000000000000000101111111111111111111111111111111111111111111111111101010000000000000000111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011001111111111111111111111111111111111111111111111111111111111111111111111110101111111111111101100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010101101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101011111111101001111111011010111111110110111111111110001001111111111101110111111101100111111101101001111111101001111111011001111111110101111111111111111101111000011110101111111110000111111101001011111111101011111111010111111111111111110111111111111110111111110100011111111110100111111101100111111111010111111111110111111111111111111001111101000000111111111000011111110110101111111101011111111111011111111111111111111000101111011001111111110010111111111000010100000000001001111111111111111111111111111111111111110100000011111111000000011111111111111111111110000000000000000000000000111111010000000000000000101101010101010101100000000000000000000000111111111111111111111111111111111111000000001111111111111111111111111111111111011111111111111111111111110101000000000000000000101111111111111100000000001101011000000000000000000000000000001011111111111111111111110101111111111111111111111111010000000000000000001011111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111011101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101111111111111111111111111111111111111111111111111111111111111111101100111111111111111010100000010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101010100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010011111111111111111010101111111111010111111111000011111010000101111111110011111111111011111111111111111010111111111011001111111010001111111111010111111110110011111010000111111111111111111111111111101010111111111101001111111100001111111011001111111110101111111111111111111111111111110011111111110100111111101001011111111101011111111010101111111111111010000011111111101011111110110011111111110001111111110100111111101100111111110001011111111111111110111111111110110111111100000000010011111111111111111111111111111111111111000001001111111000000000111111111111111111111100000000000000000000000111111111000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000101010101010101111111111111111111000001111111111111110101010000000000000000000010111111111111111100000000000100000000000000000000000000001011111111111111111111111111110000011111111111111111010100000000000000000000001111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010111111111111111111111111111111111111111111111111111111111111111011011111111111111111101100000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101001011111111100111111111110111111111111111110101111101100010111111110100101111111110100111111101100111111111010111111111111111110111111111111001111111111010011101100000101111111110101111111101011111111111111111010111111111010111111111010001111111011000111111111010011111110101011111111101111111011111111101010111111111101011111111100001111111010001011000101001111111111101111111111111111101011111111101100111111101101011111111100010011111011001111111110101111111111111110110000000001001111111111111111111111111111111111000001011111111000000001111111111111111111111111000000000000000000000111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000101111111111111110000000010101010101010000000000000000000000001011111111111111111100000000000000000000000000000000000000111111111111111111111111111111010000000101010101010100000000000000000000000010111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101011111111111111111111111111111111111111111111111111111111111111001111111111111111111010100000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000111101100111111101100011111111101001111111011001111111111000101111111111111111011111111101101111111101000111111101101011111111101001111111110101111111110111111101111110001001111111111110101111111110000111111101100111111111010111111111110111111111111111110101111111111010011111110100101111111110101111111101011111111111111111111111111111010111111111011001110100000000111111111010011111110110011111111101011111111111111111010111111111101000100111100001111111011010111111111010111101100000000010011111111111111111111111111111010000000111111111000000001111111111111111111111111110000000000000000000111111111101000000000000000000000000000000000000000000000010111111111111111111111111111111111111010110000000000000000000000000011111111111111100000000000000000000000000000000000000000000101111111111111111111100000000000000000000000000000000101111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111110110011111111111111111111101011000000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111010111111111011001111111010010111101100000111111110110011111111101011111111111111101011111111111100111111111101011111111010001111111111010111111110100101111111101111101111111111101011111111101000111111111001011111111101001111111010101111111110111111101111111111101011111111110101111111110000111111101001011111101011011111111110111111111111101000001111111110110011111110100101111111110101111111101100111111111011111111101101011110111111111111001111111111000111111111000000000001011111111111111111111111111010000000111111111000000000111111111111111111111111111100000000000000000111111111111010000000000000000000000000000000000000000001111111111111111111111111111111101100110000000000000000000000000000000011111111111111111000000000000000000000000000000000000001010111111111111111111111100000000000000000000000000001011111111111111111111111111111111111111110000000000000000000000000000000000000000101111111111111111111111111111111111100000000000101111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111110101000000000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000101000000111111101100111111111010111111111111111110111110110101001011111110100111111110110101111111110101111111101011111111111111111010111111111011001111111011010111111110000011111110110011111111101011111111101111111111111111101010111111111101001111111010010111111111010111111110110111111111101111111111111111101011111111101100111111111001011111111100001111111011010100010110111111111111111111101111111111110101111111110000111111101001011111111000010111111010111111111111111111101111111111110100000000010011111111111111111111111100000101111111111000000001111111111111111111111111111111000000000000000111111111111111000000000000000000000000000000000000010111111111111111111111111111111110100000000000000000000000000000000000000011111111111111101000000000000000000000000000000000010101111111111111111111111111100000000000000000000000010111111111111111111111111111111111111111111110000000000000000000000000000000000001011111111111111111111111111111111111111110000000000101111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111110110000000000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101101111111101000111111111001011111111011011111111100010111111111111110111111111111110011111111110100111111101000111111101101011111111010101111111111111111101111111010000011111110100011111110100100111111110100111111101101111111111110111110111111111110111111111011010111111111000011111110100011111111110011111111111011111011111111111010111111111011011111111010010010000010010111111110110011111111101011111111111111111011111111101100111111111100000100111100001111111011010111111110101111111110100000000000111111111111111111101100000101111111111000000001111111111111111111111111111111110000000000000111111111111111101100000000000000000000000000000101111111111111111111111111111111111111000000000000000000000000000000000001011111111111111111111100000000000000000000000000000101011111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000010111111111111111111111111111111111111111111111000000010111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111010110000000000000101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010110000000000000000010101001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100101011111111111111111011111111111100111111111100001111110000010111111111010111111110101111111111111111101011111111101100111111101000111111111100011111111010001111111110101100010111111111111111111111101011111111110100111111101000111111101101011111111011011111111110111111111111111110101111111110110011111110110001111111110100111111101100111111111011111110111111111010111111000101010111111111000111111110100101111111110101111111101011111111111111111111111100011011011111111010001111111111000011111110100000000000010111111111111111101000000011111111111010000101111111111111111111111111111111111101000001001111111111111111111111010100000000000000000101011111111111111111111111111111111111111110000000000000000000000000010101010111111111111111111111111011000000000000000000000001010111111111111111111111111111111111100000000000000000010111111111111111111111111111111111111111111111111111110000000000000000000000000101111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111101010110000000000000100010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101000000000000000000000010101011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100101111111110100111111101011111111111111111011111011010011001111111111010111111111000111111110100011111111101011111111111111111110111111101001001111111011001111111010000001011111010011111110110011111111111111111011111111101010111111111101011111111101001111111100001111111111001111111110101111111111111111101011111111101101111111101000111111101001011111111101011111111011000000111111111110101111111110110011111111110101111111110100111111101100111111111100010011111111111111101111111111001111111110100010100000000101111111111111110000010011111111111110110111111111111111111111111111111111111111101101111111111111111111111111111111010011001100101111111111111111111111111111111111111111111111000000000000000100110010111111111111111111111111111111111111110000000000000101001101111111111111111111111111111111111111110000000000000100111111111111111111111111111111111111111111111111111111111100000000000000010011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111010110000000000000000000100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010100000000000000000001000000000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000101111110110011111111110100111111101001011111111101011111101100001111111111111110111111111110110111111110100011111111100100111111101000111111111011010101111111111010111111111111000000111111010111111111000011111110100101111111101101111111111011111111111111111010111111111011001111111010010111111111010011111110110011111111101111111011111111111011111111111100111111111101001111111010000001011111010111111110101111111111111111101111111111101101111111101000111111101100010101111101001111111110101111111111111111111111101100000001011111111110100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000100110111111111111111111111111111111111111111111111111100101100110111111111111111111111111111111111111111111111111100000001001111111111111111111111111111111111111111111111111111111111111110110010110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101011111111111111111111111111111111111111111111111101101000000000000000101010010111111111111111111111111111111111111111111111111111111111111111111111111111010110101000000000000000001010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010011101011111111111111101011111111101101111111101001011111010000001111111011010111111110101111111111111111111111111111101011111111110100111111110000001111111101011111111011011110100000111111111111111111101111111111110011111111110100111111101000111111101100111111111011111111111111111110111111111110110111111110100011111110100101111111110101111111111011111111111111111110111111111011010000001110010111111111000011111110110011111111101011111111111111111111111111111100111101001100001111111010010111111111000111111110110010000000010111111111000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111110111101010000000000000001000101001011111111111111111111111111111111111111111111111111111010101101010000000000000000010001010011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101111000011111110110011111111101011111111111111111111111010001011011111111010001111111011010111111111010011111110110011111111111111111011111010010100111111111101001111111100001111000000010111111110110111111111111111111011111111101011111111101100111111101101011111111101001111111011001111111110111111101111111111101111111111110011111111110001111111110000111111101101011111111010111111101000001111101111111110101011111110100011111110100101111111110100111111101010111111111111010011111111111111011111111111010111111111000011110000000101111111000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000111111111111111111111111111111111111111111111111111111111010110000000000000000000001000101001010101111111111101010101010101101010100000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000001011111110110011111110100101111111110001111111101100111111110001011111111111111111111111111111001111111111010011111110100011111111100101111110100001001011111111111110111111111110111010010011001111111110010111111111000011111111110011111111111011111111111111111010111111111101011111111010001111111010010111111111010111111110101111111111111111101111111111101101111111101001011111111100011111111100000111111110101111111111111111111111111111101011111111110100111111101000111111111101010100111010111111111111111111111111111110101111101100000001011010000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111111111111111111111111111111111111111111111111111111101010110100000000000000000000000000000101010001010100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100111110101111111111111111111111111111101011111111110000111111000001011111111101011111111010111111111111111111111111111110101011111111110101101000000000111111101000111111111010111111111100001111111111111110101111111110110011111110100101111111110101111111101100111111111011111111111111111010111111111111001111111111010111111111000011111110110011111111101011111111111111111111111111111011011111111010000011111010010111111111010011111111101011111111111111111111111111111010111111101101011101001100001111111011010111111010101111111110111111000000001000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111011010101000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111010000011111111010011111111101011111111111111111111111101001100111111111101001111111100001111111111010111111110110111111111111111111011000001001011111111101100111111111000011111101000001111111011001111111111101111111111111111101111111111110101111111110000111111101001011111111101011111111110111111111111111110111111111110110111111110100101111111110001111111101100111111111010111111111110111010000101111110101111111111010111111111000011111110110101111111101011111111111011111111111110101010111111111011001111111110000011111111000011101000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000111111111111111111111111111111111111111111111111111111111111111110111111111110101011010100000000000000000000000100000001010010110100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000001010111111111001111111111000011111110100101111111110100111110110000111111111111111111111111111110101111111110001111111111000011111110100011101000000101111111101011111111111111111010111111110001001111111010010111111110010111111110110011111111101111111111111111111011111111101010111111101101011111111100001111111011001111111110101111111111111111111111111111101011111111110000111111101001011111111101001110100000101111111111111111101111111110101011111110110101111111110001111111101000111111101011001011111111111111111111111110111111111110110011111011000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111010110001010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100010111111111111111111111111111111111111111111111111111111111111010110101010010110101001100000001010101000100101101010010110100000000010101000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111011001111111111101111111111111111110111111111110101111011000000111111101101011111111010111111111110111111111111111110101111111111000010100001000101111111110100111111101100111111111010100001011111111110111111111111001111111111000011111110110101111111110101111111101011111111111111111110111111111011011111111010010111111110000111111110110011111111110011111111111011111111111111101010111111111101011110100000001111111011010111111110101111111111111111111111111111101011111111110100111111101001011111111100011111111011001111111110111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110110101010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000011111111111111111111111111111111111111111111111111111111111111111100000101010001010011010001010100000101000001001100000000000100101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111010010111111111010111111110101111111111111111111111101100101011111111101101011111111100001111111010001111111111001111111110110000000011000011101011111111110101111111101001011110110000010100111011001111111110111111111111111111111111111110110011111111110101111111110000111111101100111111111010111111111111111111111111111110101111111111000011111110100011111110110101111111101010111111111111111110111111110000011111111011001111111111000111111111000011111111110011111111101111111111111111111010111111111011001111111010010111111011010011111110110011000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111110110101010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001011111111111111111111111111111111111111111111111111111111110111011010011010001010011010100101101010010110000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111111011011111111011010011111111000011111110100101111110100100111111101111111111111111111010111111111011001111111010010111101100000000000000000011111111101011111111111111101011111011010100000011111100011111111010001111111011010111111110101111111111111111101011111111101010111111101101011111111001011111111101001111111110101111111111101111111111111110110011111111110101111111110000111111101001011111111101010000011110111111111111111110101111111110110011111110100101111111110100111111101101111111111011111111111111111110111111111111010111111111000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111101101010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001001111111111111111111111111111111111111111111111101010101010101010111010101010101010101100010100010100000000000001000000000001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100111011011111111110111111101111111110101111111110110011111011000101111111110000111111111100111111111011111111111111111110101011000000000100000001000011111111110101111111110101111110110000111010000011111111111111111011001111111111010111111111010011111110110011111111101011111111111111111011111111111010111111111100011111111010010111111111010111111110101111111111111111111011111111101011111111101100111111111001001000010100001111111011001111111110101111111111111111101111111111110101111111110000111111101001011111111011011111111110101111111111111111101000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101011010100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111010101010101010111011101010101100101010101010110100010000000100010100000000000100010100110000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000001011111100001111111010001111111110101111111111101111111111101101001011111111101101111111101001011111111101001111111011011110110000000001011010010011101011111110110101111111110000111011000000111010000101011111111010111111111111111110111111111110110111111110100011111110110001111111110100111111111010111111111011111111111111111010101111111111010111111111000011111110100011111111101011111111111011111111111111111010111100010011001111111010010111111111010111111110110111111110101111111111111111111011111111111100111111111100011111111010010111111111010111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1001010111111111111111111111111111111101011010101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111110101010010111111101010110010110011001101000000000000000001010000010000000001001010110000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100111111111011011111111010001111111010010011111111010011111111000101111111101111111111111111101011111111111101011111111010010100000000010111101100010111111111101111111111111111101111110001001011111100010001011111111100001111111011001111111010101111111111111111101111111111101011111111110100111111101000111111101101011111111010101111111110111110111111111110101011111111000011111111100101111111110100111111101100111111111100000011111111111110101111111111010111111111000011111110100101111111110101111111101011111111111111111011111111111011001111111011010110110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101101010010111111111111111111111111111111111011010101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111101101001011101011010101001100101110101010000001000000000100110000000101010100010101000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010011101100111111111010111111111111111110101111111111010111111101000011111111110100111111101101111111111011111111111111111010000000010010111110100000010110111110100011111110110101111010000101111111101000001111111111111011011111111010001111111010010111111111010011111110101011111111111011111111111111101100111111111101011111111100001111111011001111111110101111111111101100111111111111101011111111110100111111101000111111101100000011111011011111111110111111111111111111101111111110110011111111110001111111101000111111101100111111111010111111111110111110111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111110101011010010101111111111111111111111111111111010110101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010011111111111111111111111111111110101101010101001010101111111010110101001011000000000101000100010010110101010000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111101001011111111101001111111011001111111110111111111111110100101111111111110101111111110000111111101000111111111101010000000000111111111011000100101111111110110111111110110101101000010011111111110001011111111010111111111111111110111111111110101111111111010111111110100011111110110101111111101010111111111011111110111111111010111111111010001111111010010111111111000101111110110011111111101011111111111111111010111111111100000101111100001111111010001111111111010111111110101111111111111111101011111111101100111111101001011111111100011111111011001111111010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111010110100101011111111111111111111111111111010110101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000111111111111111111111111111111010010111111111111111111101101010100101100000000000001001010100100110101010000010100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111111010111111101101011111111100001111111111010111111111000011111111101111111111111111111011111111101100111111101100000001010111111111111100000111111110101111111111111111101110100100101111111111100000111111101001011111111101001111111010101111111110111111101111111110101011111111100101111111110001111111101000111111111010111111111010111111111111111110101111111111000111111110100011111110110101111111110101111111111010111110100000111011111111111011001111111010010111111111000011111110110011111111101011111111111111111011111111111011011111111100001111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111101110110101001010111111111111111111111111111110101101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000001111111111111111111111111111101111111111101110111011000101010001000000000000010101010011000100101100000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001011101100111111111010111111111111111110111111111111001111101100010111111111000011111111110011111111101011111111111110110000000100111111111111110000001111111111000111111110110011111100000101111111111111000100111111111010111111111101011111111010001111111011010111111110110111111111101111111111111111101011111111101100111111101001011111111101001111111011001111111110111111010111111111101011111111110101111111110100111111101000111110100001011111111010111111111111111110111111111110110111111110100101111110110001111111101000111111111010111111111110111111101111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111010101101001010111111111111111111111111111110101100110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000011111111111111111111111010101010101101010001010101010000000000010000000000010101001010110100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100101111110000111111101001011111111101011111111010111111111111101100101111111110110111111110110101111111110000111111101100000001001111111111111110100100111111111111001111111110100011110100010011111111111111000011101010111111111111111110111111111010101111111011010111111111000111111110100011111111110011111111101111111111111111111010111111111101011111111010001111111010010101011111010111111111101111101111111111101011111111101100111111110000011111111101001111111011001111111110101111111111111111111111111111110011111111110100111111101001011111111101001111111010100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111110101100110010101111111111111111111111111110101011010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000001011111111111101011010100010000000001010100101010111011000000010101000001001011111110101000000000000001010100000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111010111111101100111111111101001111111010001111111011000111111110101111111111111111101011111111101101111111000000000011111111111111111011000011111111011111111111111110111111000100101111111111111110010111110000111111101001011111111010111111111111111110111111111110101111111110110011111110110101111111110100111111101100111111111011111111111111111110101111111111000000111111010011111111000011111111110011111111101011111111111111101001001111111011011111111010001111111010010111111111010011111111101011111111111111111011111111111100111111111101001111111010000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111110111011001100101111111111111111111111111111111011010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111101000000010000000001010101010101010101000000000000000001010010110100000000010101000100111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100111110110100111111101011111111111111111010111111111011011111111100010111111111000011111110110011111111101011111111110100000001011111111111111111111100001111111010010111111111010111111100000111111111111111111010010111101011111111101100111111111100011111111100001111111111001111111111101111111111111111101011111111110101111111110000111111101001011111111101011111111110111111110000111110101111111111110011111110100101111111110001111111101100101000010010111111111111111110111111111110110111111111000111111110100101111111110101111111101011111111111111111110111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111101010110101001011111111111111111111111111111010110100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111111111110110100110010101011001100110011010001010101010000000000000000010000000001010000010111101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010010111111100101111111110000111111101101011111111010111111111111101010111111111110101111111110100011111110100101111011000000001011111111111111111111101000001111111010111111111111010111101000010011111111111111111100000011111111111111111111111111111010111111111011001111111010010111111111010111111110110011111111101111111111111111111011111111101100111111111101011111111100001111110001001111111110101111111111111111101111111111101011111111101000111100000001011111111101011111111110101111111111111111111111111110110111111110100101111111110000111111101101011111111100110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111010101101010010111111111111111111111111111110101101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001001111111111111111111111111111111110101100101111111111110000000000000001010000010100010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100101111111111101011111111101100111111101101011111111101001111111011001111111110111111101111111111101111111111110010110000000100111111111111111111111110100101111010111111111110111110111110100100111111111111111111111100000100111111110000111111101010111111111110111111111111111110101111111110110111111111010011111110110101111111110101111111111011111111111111111010111111111011001110100000010111111111010111111110110011111111101011111111111111111011111010000100111111111101001111111100001111111011010111111110101111111111111111111111111111101010111111101100111111111100000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111110101100101010111111111111111111111111111110101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111110101010101111111011010100010000010101001011000000010101010100110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101111110100011111111101011111111111111111011111111111100111111111100001111111010010111111111010111111111101111111101000000001111111111111111111111111111000101111100001111111011010111111010010011111111111111111111101001001011111111101101111111101001011111111001011111111011011111111110111111111111111111101111111110110011111111110101111111110000111111101100111111111010111111111111000010111111111110110111111110100011111110100101111111110100111111101100000101111011111110111111111110101111111110001111111111000111111110100011111111110011111111111011111110111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110101011010100101111111111111111111111111111101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000001010111111111111010110101010010101010101100000000010101001011101011000001001010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001010111111111000011111110100101111111111111111111111010111111111111101010111111111110101111111111010011111111000100110000000101111111111111111111111111111010010111111010111111111011001111101100010111111111111111111111101001011111101111111111111111111011111111111011011111111100001111111010001111111111010111111110101111111111111111101011111111101010111111101000111111111001011111111010010111111110101111111111101111101111111111101011111111110001111111110000000001101101011111111010111111111111111111101111111110101011111110110011111110100100111111110100111111101100111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111101010110100101011111111111111111111111110101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000100111110110100010001010100000000010000010001000100000000000000000001010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111110111111101111111111101101111111111111111111101001011111111101001111111010101111111110111111111111111110100000000001001111111111111111111111111111111100001100111111111110111111111110110000101111111111111111111111110100111110110101111111101101111111111011111111111111111110111111111111001111111011010111111111010011111110110011111111101011111011111111111111111111111011011111111100001111111010001111111111010111111110101111111111111111111111111111101010100000111000111111111100011011111101001111111110101111111111101111111111111111101011111111101100111111101000010000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101001011111111111111111111111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000010010110011101111101100000001001111111111101011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010011111110110011111111111111111111111111101010111111101101011111111100001111111011010111111110101010100000010011111111111111111111111111111111110001001001011111111101001111111011000011111111111111111111111111110001111111110101111111110000111111101000111111111101011111111110111111111111111111101111111110110011111110100101111111100101111111101100111111101010111111111111101000001111111011001111111111010111111111000011111110110101111111101011111111110001011111111111111010111111111010001111111010010111111111010011111110110011111111101111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000100010101001011000100101000001111111010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011010111111111000011111111000101111111111111111111101011111111111111101100111111111010111111111011010111111110000000000100111111111111111111111111111111111110110001111011111111111101011111111000001111111111111111111111111111100000101111111111111111111111111111111100111111101101011111111100001111111011001111111110101111111111111111111111111111101101111111110001111111101000111111111100001001011010111111111111111110111111111111101111111110100011111111100001111111110001011111111100111111111011111111111111111110111111111111010111111110100011111111110101111111101100111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000101000001000101010000000101000001010011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011010010111111111111111111101011111111111111111111110000111111101001001111111010111111111111101111111111111011000000001111111111111111111111111111111111111110100001111111111011111111111110110001011111111111111111111111111110110001000011111111110101111111101110111111111111111011111111111010101111111011010111111110010111111111010011111111101011111111111011111111111111111100111111101100000000111100001111111011010111111110101111111111101111111111111111101011111111110000001111101001011111111101001111111011011111111110111111111111111110101111111110110101111111110001010000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000101001110101100000000000000000001010100000000000000000000000000010010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010101011011010111111110110111111111111111111111111111101011111111101001011111111001001111111101001111111111001100000101111111111111111111111111111111111111111010000000111111101001011111111011000101111111111111111111111111111110100100110011111110100101111111110101111111101100111111111010111111111111111110111111111110101111111111010011111110100101111111110101111111101010111111111111111110100000111010111111111010001111111110010111111111010011111111110011111111111011111000001111111010111111111101011111111100001111111010001111111011010111111111101111111111111111101000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000001110110100000001001011000000000000000000000000000000000100111010110000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001001011000100111011010111111011000111111110100011111111110011111111101111111011111111111010111111111101001111111100000000001111111111111111111111111111111111111111111100001011111111101100111111111000010011111111111111111111111111111110100101111111101111111111111111101100111111101000111111101101011111111011001111111111011111111110111111111111111110110111111110110101111111110000111111101000111111000000111111111010111111111111111110101111111111010011111110100011111111100101111100000100111111111011111111111111111110111111111011001111111111010011111111000011111110110101101000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000001001100010100000100000000010100000001000000101110110000000001001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111010100111111111111111110101011111110110011111110110101111111110100111111101100111111111011111111111111101100000100111111111111111111111111111111111111111111101001011111101011111111111111101001001111111111111111111111111111111111000101111110110011111111101011111111111111111111111111111010111111111101001111111010001111111011010111111110101111111111101111111011111111101011111111101101011110000001011111111101001111111011011111111110101111111111111111101011111110110101111010000000111111101000111111101101011111111010111111111111111110101111111110110011111110100001000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111111111101000000000000001001100000001010100000100111110110000000001001100000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100001101011010001111111011001111111110111011111111111111101011111111110100111111110000111111111101011111111011000000001111111111111111111111111111111111111111111111110000111111110000111111101101000000111111111111111111111111111111111111000101111110100011111110100101111111110101111111101010111111111011111110111111111010101111111011010111111111000011111110110101111111110011111111101011111111111010010010111111111011011111111010010111111011010111111110110011111111101111111111111010000101111111101100111111111101011111111100001111111011001111111110101111111111111111110000000000000101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000001010011111111111111111111111111111011110100000000000000000101010100010100111011010000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101011010100111101001111111010010111111111010111111110110111111111101111111111111111111011111111101101011111101000000101111111111111111111111111111111111111111111111110100101111111101101111111101000000111111111111111111111111111111111111111000101111110111111111111101011111111110000111111101000111111101101011111111010111111111110111111111111111110101111111110110011111110110101111111110100111111101100010111111011111110111111111110111111111111010111111111000011111110100101111111110000000011101011111111111111101010111111111011011111111010010111111011010111111110110011000000000000000000000101010101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000101001111111111101111111111111111111010110100000000010101000001000001000100000000000000010100101100000000000011010000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000111111000100111110111111111110101111111111010111111111000011111110110101111111110010111111111011111111111110100000001111111111111111111111111111111111111111111111111111000011101011111111111111111100010111111111111111111111111111111111111111000101010111111110101011111111101111111111111111101010111111111000101111111100001111111010001111111111001111111111101111111111111111101011111111110101111111101000001111101101011111111011011111111010111111111111111110101111111110110011111110100100000101110000111111101100111111111010111111111111111110111111111111010111111111000010100000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000101010011010001001111111111111111111111101101010010000000000000000000000000000000111111110000000100010011000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101001001101001101001111111011001111111110111111111111111111101111111111110011111111110100111111110000111111111100000101111111111111111111111111111111111111111111111111111100010111100101111111110100110000011111111111111111111111111111111111111111000001000111111110100011111110110101111111101011111111111011111111111111111010111111111011001111111010010111111111010011111110110011111111101111111111111111101001011111111101011111111100011111111010010111111111001111111110101111111111111111101010100001101101111111101000111111101001001111111101001111111110101111111111111111101111110000010001000000000000000000000000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101000000000000000000000100101010101010101011010101010000000000010101000000000000001101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101010110100101101011111111100001111111010010111111111010111111111101111111111111111101011111111101100111110110000001111111111111111111111111111111111111111111111111111111001001111101101111111110000000100111111111111111111111111111111111111111111000100111111111110101011111111110011111111110001111111101000111111101100111111111110111110111111111110101111111111010111111111000011111110100101111111110101110001001011111111111111111011111111111011001111111010010111111111000111111110110011111111100001111111111111111011111111111010111111111101011111111010010111111111010011111110110100101110110010101010110011010000000000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101001110101101000000000000000001000000000000000000000001010100101111010000000001010100000000000000000000010100010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100110100111111000001111111111111111010111111111010101111111111010111111111000011111110110101111111101011111111111011000000111111111111111111111111111111111111111111111111111111101000001011111111111111111100000011111111111111111111111111111111111111111111000101111110101111111111101111101111111111101011111111101100111111101001011111111100011111111011001111111110111111111111111111101111111110110011111111110000110000101000111111101101011111111010111111111111111110101111111110101011111110100011111110100000111111110100111111111010111111111111111110111111111011001111111010010111111111000000111111100101111111101101101110100000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000010011111010010001001010101010000000000000000000000100101010110001001010101010000000000001001100000000000100000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000111100010001011111101101011111111010111111111111111011101111111110110111111110110101111111110001111111110000010111111111111111111111111111111111111111111111111111111110100101000011111111110101101100010111111111111111111111111111111111111111111111000101111011000111111111010011111110110011111111101111111011111111111011111111111100111111111100001111111010010111111111010111111111101111111111111111101110100001101100111111101101011111111100011111111011001111111110101111111111111111101111111111110001011111110100111111110000111111111001011111111010111111111111111111111111111110101101011110110101111111100100111010110000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000001010001011111101101001101001010101101000000000101000000001101010011010000000000101011000000010000010100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100101111101011110000101100111111101001001111111100001111111011001111111110101111111111111111101111111111110010111111000000111111111111111111111111111111111111111111111111111111111110100011110011111110110101110001001111111111111111111111111111111111111111111111000101111110101111111110110011111110100011111110110100111111101100111111111011111111111111111110111111111111001111111111010111111111000011111110110011111111000101111111111111111011111111111100111111111100001111111010010111111111010011111110101011101000001111111011111111111010111111101100111111111100001111111010001111111111001111111111001111111111111111110101111010101100111101000000000101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000001010101001010101111101011010001000101010011010000010100000000000000000100110100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001011110101111111000101111111111111111011111111111010111111111010001111111110010111111110110011111111101011111111111100010011111111111111111111111111111111111111111111111111111111111110000011111111111111111110100101111111111111111111111111111111111111111111111110100001001111111110101111111111111111101011111111110101111111110000111111101001011111111101011111111110111111111111111110101111111110101011111111100101111111000100111111101100111111111010111111111111111111111111111110101111111111010111111110100011111000000101111111101011111111111111111110111111111010111111111011010111111010010111111111000011111110110011110011111101011011111110101000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001000001001110101101010100101001001111101101010001010000000000000000000000000000010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100111110100101101100000000111111101000111111111100111111111111111111111111111110101111111111010111111110100101111110110001011111111111111111111111111111111111111111111111111111111111111010010111111110100011111010000011111111111111111111111111111111111111111111111111000000010111111111010111111110110111111111101111111111111111111011111111111100111111101101001111111100001111111111001111111110101111111111111111111111111010000101111111110000111111101000111111101101001111111010101111111110111111101111111110110011111100000101111111110001111111110000111111111100111111111011111111111111111110101111111111000011111110100101110101100000011111101101111011000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0000101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000100000001001111101100010100010000101111100000000001001101000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001011111111111011110101110101111111101000111111101101011111101101001111111010101111111110111111101111111110110011111010000101111111111111111111111111111111111111111111111111111111111111111100001111111110110011111010000101111111111111111111111111111111111111111111111110100100111111111011010111111111000011111110100101111111110101111111111011111111111111111110111111111010101111111010001111111111010011111110110011111110101100010111111111111111111111111100111111111101011111111100001111111011010111111110101111111111111100010111111111101011111111101100111111101101011111111100011111111011011111111110111110110111111111101111110100101101011111110000111111101000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0110100000101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000001001101000101001011000100010101000000000000010100000000000100101100000000010100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100111111000011111111000101111111111011111111111111111010111111111101011111111010001111111111010111111110101111111111101001001111111111111111111111111111111111111111111111111111111111111111101101011110111111111111101100001111111111111111111111111111111111111111111111111111000101111110111111111111111111111111111111110011111110110101111111110000111111101100111111111010111111111111111111111111111111001111111111000111111110100000010111110100111111101011111111111111111110111111111010101111111011001111111110010011111111000000000111110011111111101111111111111111111010111111111100111111111100001111111010010110110010110111111111110000111011001111111011111111101101000000000101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111101010110101010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100000000000001010100101101010000000000000001000000000000000101000000000001001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011111110110011111100000101111111110100111111101100111111111110111111111111111010101111111111010111111111000011111110100000111111111111111111111111111111111111111111111111111111111111111111110000111111010011111110110000111111111111111111111111111111111111111111111111111110100001111010001111111111010111111111111111111111111111111111111111101011111111101000111111101001011111111011001111111110101111111111111111111111111111110000001110110101111111110000111111101000111111111010111111111111111111111111111110101111111110110100000110100101111111110101111111101101111111111011111111111111111110111111111111001111110101000011111110100000111111010101111111101011111111101000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111011010101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010101010000000000000000000000000100110011010000000000000000000101010100000000000101010000000000000000000100000000000000000100000000000000000000000000000000000000010100101110101111101111110100101011111110110100111111110000111111101101011111111100111111111110111111111111111110101111111010000111111111111111111111111111111111111111111111111111111111111111111111110101111111010111111110100100111111111111111111111111111111111111111111111111111110110000111011001111111011010111111110111111111110110011111111101011111111111111111111111111111010111111111101001111111010001111111111010111111110101011101000001111101111111111101011111111101100111111101100011111111100001111111111001111111110111111111010000011101111111111110101111111110000111111101000111111111101011111111110111111111111110101101111111110110001011111000001111111110000111111101000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101011001100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101000001010101010101010101010010101010000100000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000001000000010011111111010011111111000101111111101111111011111111111011111111111101011110111100001111111010001111111111001111111111110001001111111111111111111111111111111111111111111111111111111111111111111110100010111111111111111011000011111111111111111111111111111111111111111111111111111111100000111111111111111111111111111110111111111110100011111110100101111111101001111111101010111111111011111110111111111110101111111011010011111111000011101000000011111111110011111111101111111111111111111010111111111011001111111010010111111111010011111110000011111111101111111111111111111011111111101100111111101100011111111100001111111111000000111110101111111010001110100111111111101101111111101100101000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101111111111111111111111111111111111111010101011001011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000101111111101100110100000000010000000000010100000000000000000000010100000000000000000000000000000000000000000000000000000000000000000100000000000101001111111011010011111010000011111110100101111111110010111111111011111111111100111010111111111011001111111010010111111011000101111111111111111111111111111111111111111111111111111111111111111111111010001010010111111111010100010111111111111111111111111111111111111111111111111111111111110000011111111011001111111110101111111111111111111111111111101011111111110100111111101000111111101101011111111011011111111111111111111111111110101111110000010011111110110100111111110001111111101100111111111011111111111111111110111111111011010111111111000011111110100011111111110101111111111011111111111111111110111111111011001111111010010100111111000011111011000101110011101011111111111111111011111011000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010100101011111111111111111111111111111111111111111010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000101001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111110101111111111101001001011111110110101111111110001111111101000111111110000111111111110111111111111111110101111111100010111111111111111111111111111111111111111111111111111111111111111111111111010001011001111111111000001001111111111111111111111111111111111111111111111111111111111110001011111111010001111111010010111111111111111111110101011111111101111111111111111111010111111111101011111111101001111111010001111111111001111111110110000111111111111101011111111101100111111101000111111101101001111111011011111111110101111111111111111000101111110110011111110110100111111110000111111101101011111111010111111111110111111101101011111001111111111000011100011100101111111110100111111111100110000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1001101010101010010101011111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000010100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100001111111100010111111111000100111111101111111111111111101011111111101100111110110001011111111101001111111011001111111110110001001111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111110100000111111111111111111111111111111111111111111111111111111111111110001011011111111111111111110101111111110111111111110100011111111101101111111101101111111111011111111111111111010111111111011001111111011010011111111000000111110110011111111101111111111111111111010111111111101011111111100011111111010001111111111010110100000101111111111111111101111111111101101111111101001011111111100011111111011001111111011001111111110111111000011110011110011111111110100111111101001011010000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111101011010101000101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000010011101010101010110101010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000010010111110101101001111111010000011111111000011111110110011111111101011111111111011001110111111111101011111111010001111111011000100111111111111111111111111111111111111111111111111111111111111111111111111101000001111111011001111000101111111111111111111111111111111111111111111111111111111111111110001001101001111111010111111111110111111111111111110101011111111111011111111110100111111101000111111111100111111111010111111111111111110101111111111000000111110100011111110100100111111101101111111101011111111111111111010111111111011001111111111010110100000000011111110110011111111101011111111111011111111111111111100111111111100001111111010010111111111010110110011100101111111111011111111111111101100111110110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111101010110101010100101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000000100101111111111111010110000000000000000000000000000010100000000000000000000000000000001000000000000000000000000000000000001011011111011010011111111101100001111111110110011111110100101111111110101111111101000111111111011111111111111111010111111101100010111111111111111111111111111111111111111111111111111111111111111111111111111101001011111111010001010010011111111111111111111111111111111111111111111111111111111111111101000011101011111111100001111111010111111111110101011111111111111111111111111101011111111101100111111101101011111111100011111111011001111111110111111000001011110101111111111110011111111110001111111101001011111111101011111111010111111111111111110101110100001010111111110100101111111100101111111110100111111111010111111111011111111111111111110010111111111010011100101000101111110110101111111101101111111111011101100000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101010101011001100101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101000000000100110100010100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000001010001011111101000001111111011000000111110101111111111111111101111111111110101111111110000111111101001011111111101011111111110110001011111111111111111111111111111111111111111111111111111111111111111111111111111100101111111111111101100010111111111111111111111111111111111111111111111111111111111111111101000011111111111111010111111111011011111111110110111111110101111111111110011111111101111111111111111111010111111111011011111111010001111111010010110000000010111111110101111111111111111111011111111101100111111101001011111111100001111111010001111111111000100111111111111111111111111110011111111110101111111101001011111111101011111111010101111010111111111101111110100110100111111110101111111110000111111101001011011000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111101010101011010100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000100111010111111010101001111111010000101111110010111111110110011111111101011111111111111010011111111101100111111111100011111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111000011111101001111101000001111111111111111111111111111111111111111111111111111111111111111111000001111111011011111111110111111111111111110101111111110101111111110100101111111110001111111101100111111111010111111111111111010111111111111001010000000010111111111000011111110110011111111101011111111111011111011111111111011011111111010001111111010000000111111010011111111111011111111101111111011111111101010111111111101001111111100001110100100010111111110100001111100101111101111111111101010111111101000111111110000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110101010101101001100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101100000000000000000101010000000000000000000001000000000000000000010000000000000000000000000000000000000001000000111111101101001111111110111010010111111111001111111111000111111110100011111111110101001111101011111111111111111011111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111010011111101001111100001011111111111111111111111111111111111111111111111111111111111111111111100010111101100011111111101001111111111001111111110101111111111111111101111111110101010111111110000111111101001011111111101011111111010111111111100000001001111111110110111111110110101111111110001111111101100111111111010111111111111111011101111111110100000111111010111111111101011111110110101111111101101111111111011111111111111111010101111110101001111111110000000111100010011111110110011111111101011111111111111110000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111101110101010110010110010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100000000000001001100000000000000000000000000000000000000000000000000010000000000000000010000000100110100111111010000011111111101001000001110101111111111111111101111111110101011111111100000111111110000111111101100111111111010110000111111111111111111111111111111111111111111111111111111111111111111111111111111111010101111111110111111000100111111111111111111111111111111111111111111111111111111111111111111111100010111111010111111111011001111111010010111111111010111111110111111111111101111111111111111111011111111111100111111111101001111111100001111111100000001011110101111111111111111101111111111110011111111110000111111101001011111111101001111111011011111110001001111101111111111111011111111110101111111110000111111101101011111111100111111111110110101111111111110101001011010010011111110100101111111100100111111101101010000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111010111011010101001010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101100000000000100000000000000000000000000000000000000000000000000000000000000000000000001001011101011101101001100111111111100000001011010010111111111010111111110101111111111101111110101111111101101111111101000111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111011001101011111111010000111111111111111111111111111111111111111111111111111111111111111111111111100010100111111111011111111111111111111111111111011010111111110111111111110100101111111110100111111101011111111111111111010111111111010101111111100000001011110010111111111010011111111110111111111111111111111111111111100111111111101011111111010001111110000010111111110110111111111101111101111111111101011111111101100111111101100011111111100000101111011001111111100001011001111111111101011111111110101111111110000000001000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101011010100110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101000000000000000000000000000000000000010000000000000100000000000000000000010100110100111110100000111111111011111010000101111011001111111011010111111111000011111110100011010111101011111111111111111110111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001101011111111100010111111111111111111111111111111111111111111111111111111111111111111111111010000000111111111100011111111011011111111110111111111111111111111111111110110011111110110101111111110000111111111101011111111010111111111111111000010001011110110111111111000011111110100101111111110100111111101011111111111111111010111111111011011111101000010111111111000111111110110011111111110011111111111111111111111111111010111111111011001100111010010111111010000011011110110011111111101011111111111110110000000001010000000000010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011010011001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101000000000000000100000000000000000000000000000000000000000000000001001111100000111101000000111111101101011010000100111111111111111110111111111110101111111110110000001111100101111111110000111111101010110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101011011111111101001001111111111111111111111111111111111111111111111111111111111111111111111111010000101111111111100111111111100011111111010010111111111010111111110101111111111111111111011111111101011111111101000111111101100011111111101010001001000001111111111111111111111111111101011111110110101111111110000111111101000111111111010111111111110101001011111111110101111111110100011111110100011111111110011111111101100111111111011111011101101011010111111111111000110110111000011111110100101111110110101000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101100101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010110100000000000000000000000000010000000000000000000000000101101111111011110100101100111111101101001001001100001111111011001111111110101111111111111111101001011111101011111111110101111111101000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000111111111100110000111111111111111111111111111111111111111111111111111111111111111111111111111111000011101011111111111111111110111111111010101111111110010111111111000011111110110011111111101011111111111111111011111111111010111111111100000001001000010111111011010011111110101111111111111111111011111111101011111111101101011111111000011111111100010001011011001111111111111111111111111111101011111111101111111111101000111111101101011111111001011111111110111111000010110111101111111110110011111110100000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101011010100000000000000000000010000000100000000000101010101111010000101111111111011111010110000111010111111111010001111111010010111111111000111110100101011111111101111111111111111101100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111101000000000111111111111111111111111111111111111111111111111111111111111111111111111111111000011101000111111101100111111111010111111111111111111111111111110110111111110100101111110110001111111110100111111111010111111111110111111110000111000001111111111010111111111000011111110110101111111101011111111111011111111111111111011111111111011010001011010001111111011001111111110110111111111111111111111111111101011111111111101011111101100001111111010010110100101010111111110101011111111111110100000000000000000000000000000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101010101100010000000000000000000000010101000101101101000000111111110000111011000000111111111110111111111111111110111111111111010110110100100011111110110101111111110011101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111011000101111111111111111111111111111111111111111111111111111111111111111111111111111110100101101100111111111101001111111100001111111011001111111110101111111111111111111111111111101011111111110100111111101000111111101101011111110001111100010111111110111111111110101111111110110011111110100100111111110001111111101100111111111011111110111001011110101111111110101111111111000011111110100101111111101101111111111011111111111111111011010111111011011111110000000111111111000011111110100100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101101000001010101010011111011000100101101111111101100101100000001011111111101001111111010101111111110111111111111010110101111111111110101111111110001000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101101111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111100101111111111111111011111111111010111111111010001111111010010111111111010011111111110111111111111111111111111111111101111111111101011111100001111100010100001111111111001111111110111111111111111111101011111111101100111111101000111111101100011111101000011111111110111111111111111111101111111111110011111110110001111111110000111111111101011111001010111111111111101001010011111111010111111110100000000000000000000000000000000000000000000101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000010110100000100111100000011111011010010111011101000010010111111111101011111111010001111111011010111111010010111111111101111111111111111101100010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101110000111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111101100111111111010111111111111111111111111111110101111111111010011111110100101111110110101111111101101111111111011111011111111110101111010000011010111111010010111111111000011111110110011111111101111111111111111111010111111111101011111111000001111111010010111111111010111111110101111111111111111111011111111101101111111101001011110110000011111111010010001010100101111111111101110100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010001010101000000010100110001000101111010000000010010110001011111111011111111111111111010101111111111001111111100000011111111000011111111110011111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011101011111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011111101000111111101101011111111101001111111111011111111110111111111111111110101011111111100101111111110000111111101000111111111101000001111010000010111111111110111111111111010111111110100101111111110101111111101101111111111011111111111111111001011111111011001111111011010111111110100111111110110011111111101011111111111111111110111110110101011111111010001100010100000111111111000101000000000000000000000000000000000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000011010000010011111111000011110111111110110100000000000001011111101001011111111101011111111110111111111111101101001111111110110111111110100101110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111101001001111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111111111111111010111111111101011111111100001111111111010111111110110111111111101111111111111111101011111111101100111111101000000101111011000101111011001111111110111111111111111110101111111110110101111111110000111111101000111111111101011001011010111111111111111110101111111110110011111110100101111111110100111111101100111111111010110011111111111110111100010101010111111111000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000010111101100000111111111101111111011110000000001010111101100111111111100011111111100001111111011000011111110101111111111111111101111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000100111111101010111111111110111111111111111110101111111011001111111111000011111110110011111111110011111111101111111111111111111011000101111111000001111100001111111010010111111110110111111111101111111111111111101011111111101100111111101001001000111100011111111011001111111110101111111111111111101111111111110101111111110100111111101001010101111101001111111010010100111110111110110000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000010100000101001011010110110000010011111110100101111111110001010000000000101111111111111010111111111011011111111010010111111111010111111110110011111010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101111110100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111111101000111111111101011111111011011111111110111111111111111110101111111110110011111110110101111111110100111111101100111111000101111110100000111110111111111111001111111111000011111110100011111111110101111111111011111111111011111111101001011011011111111010010111111110010111111111010011111111101011111111111111111011111111111100101101111100011111111100000000111011010111000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110100000001000000001011111110111011000011110111111110100011111110100001011111000000000100101100111111111010111111111111111011001111111111010111111111000011101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101011000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010011111111101010111111101100111111101101001111111010001111111011001111111110101111111111111111101011111111110101111111101000111111000101111111100001011111111010111111111111111110101111111110110011111111100101111111110001111111101100111111101001011111111111111110111111111110101111111110100011111110100011111111110100111111111101111111101100111111111111111011000000111010010011000000000000000000000000000000000000000000000000000001000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000000100111111111111101000010111111110101111111111111110100001111111101101000000000001001111111001011111111011001011011110101111111111111111101111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011101101111111111011111111111111111010111111111011001111111010010111111111000111111110110011111111101111111111111111101011111111000101111111110000011111111100001111111011001111111110101111111111111111101111111111101101111111110000111111101001011111111101001111111010101111111110111110111111111110110011111111110101111111110000111111101001011111111101011111110001011111101000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010100110010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101000000000000000101001111111111111110110100010111111111000011111110110100000101101011111111101001000000000101001101011111111100010101111010010111111111010111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101110101111111101000111111101100111111111010111111111111111111111111111111010111111111000011111110100011111111110101111111101010000101111111101000001111111011001111111110010111111111010011111110110011111111101011111111111011111111111111101001011111111101001111111010001111111011010111111110101111111111101111101111111111101011111111101001011111111000001111110000010111101000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101010101011010010110011010010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000000000000000010101001011111111111111111111000010101111111111010111111111000000010111100101111111110000101101000000000011111110111010110101111011001111111111010111111010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000101011111111101100111111101001011111111101011111111011001111111110101111111111111111101111111111110011111111110100111111101000000011111111101000010010111111111111111110111111111111010111111110100011111110100011111111110101111111101010101000111011111110111111111011001111111111010111111111000011111110110011111111110011111111101111111011011111111010111111111000001110100000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111010101010101010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010000000101010101001010101011111111111111111111111100010111111110101111111111111110100001011111110011111110110100111110110000000000010101011110110000111111111111111110101111101001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111101011111111111111111011111111111101011111111100001111111010001111111111010111111110101111111111111111101011111111101000000011111111111010000001011111111011001111111110101111111111111110101111111111110011111111110000111111110000101000111101011111111010111111111111111110111111111110101111111110100011111111100101111111110000111011010100111111111010111100001111000000000000000000000000000000000000000000000000000000000100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000100111011111111111111111111111111111111111111110000001111111010010111111111010011000100101011111111111111111011111111101100101100000000001111000000001111111011001111111110100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111110101111111101101111111111011111111111111111110111111111011001111111011010111111111000011111110110011111111101011111011000011111111111010000001011111111100001111111010010111111111010111111111101111111111111111101111111111101011101001001001011111111100001111111100001111111110101111111111111111111011111111101011111111101100111111010001011111111001001010010010000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010100111111111111111111111111111111111111111111111111000100111111111111001111111111000100010110100011111110110101111111101011111111111011010000000100010010111111111010001111111010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111110101111111110000111111101001011111111101011111111010111111111111111110101111111110110111111111100101111111100101111110000101111111111011000001111111111110111111111111001111111111010111111111000011111110110101111111101011111111101000111111111111111010111111111011001111111010010111111011000011111110110011111111101111101111111111010010111111111101011111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101010010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000111111110111111111111111110101000001110110011111111100101111111110000111111101000111111000000010100111111111111111111111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010011111111111111111011111111101010111111111101011111111100001111111011001111111110101111111111111110111111111111101101111010000100111111111110100000111101011111111010111111111111111110101111111110110011111110110011111111100001111111110001011111111100111111111111111110111111111110101111111111010111111110100011111110110001111111101100010111111010111110111110100000000000000000000000000000000000010000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101010101101010101010101001010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111100001111111011010111110000001111111111111111111111111111110011111111101000111111101000000000010101001111111010101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111110101111111101011111111111111111011111111111010111111111010010111111011010011111110110011111111101011111111111010000011111111111110100001011101011111111100001111111011010111111110101111111111111111111011111111101011111111110000111111101001011111101100011111111011011111111110111111111111111110101011111111110101111111110001010111101001011111111100000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111101110101010110101010011001010101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011111111011011111111010001110110000000111111110100011111111101011111111111111111111111111110000101000000000001111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100111111100101111111110001111111101100111111111010111111111111111110111111111110101111111111010011111110100101111111110000000111111111111111110001011110111111111010111111111011001111111110010111111111010011111111110011111111111111101001011111111011111111111101011111111100001111111010010111111111010111111111101111101111111111101010110111101100111111101001010000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111101010101010101101010100101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000111010111111111111111111101111000001001111111111010011111110100101111111110001111111101101010111111010110000000100111010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111101101111111101001011111111001011111111101001111111110101111111111111111101111111110101011111110110000000011111111111111101000001011111010111111111111111111111111111110101111111110110011111110100101111111100100110000101101111111111011111111111111111010111111111011001111111111000011111110100011111111110011111110110101111111111111111010110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111101010101011001011010011010010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111001011111111010001111111010000011111111111111111111111111110011111111110100111111110000001111101101011110100000010100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010011111111101011111111111111111111111111111010111111111101011111111010001111111111010111111110101111111111111111101010000011111111111111101000010111101001001111111100001111111010101111111111101111101111111111101111111111110101110000110000111111101000111111111100111111111110111111111111111110101111111110110011111110100101111111110000111111101100111111101000000000000000000000000000000000000000000000000000000000000000010011111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110111011101010110011001100101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010011111010111111111101001111101000010111111111010011111110101011111111111011111111111111101001001111101101011111111000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000011111110100101111111110101111111101011111111111111111111111111111010101111111011010111111111000011111110100011111111000011111111111111111010000011111010111111111011011111111010010111111111010111111110110111111111101111111111110000101011111111101100111111101100011111111100001111111011001111111110111111111111111111101111111111110100111111110001011111110000000000000000000000000000000000000000000000000000000000000000010011111111111111111111111111111010110101001101010101000101010011010101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110110010101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100001010111111111111111110111110110001001111111111010111111110100011111110110101111111101010100001011111111011111111111011000100000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111101011111111110100111111101001011111111101011111111010111111111111111111111111111110101111111110110101111111000100111111111111111011000100111111111111111111111111111010101111111011010111111111010011111110100011111111100101111111111011111111111111111011111111111010001110101100000101111111000111111110110111111110101111101101111111111011111111101000000000000000000000000000000000000000000000010000000000000001001111111111111110101011010100000000000000000000000000000000000000000000000000010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000101000111111111101011111111011000000111111111111101111111110110111111110110011111111100000000000101000111111111100111110010111101100000100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000101011111111111111111011111111101011111111101101011111101100001111111010001111111110101111111111111111111111111111000101111111111111111111000000111111111101011111111011011111111111111111111111111110101111111110110011111110100001111111110100111111101100111111101010101011010100000001010011111111010111111111000011111110100101101101110100111111101010111100000000000000000000000000000000000000000000000000000000000000001111111111101101000000000000000000000000000000000000000000000000000000000000000001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100111100111111101001011111111100000011111010001111111110110111111111101111111111111111101001000001110100111111101001011101011111111111010000010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000011111110110101111111101011111111111011111110111111111010111111111011001111111010010111111111010011111110110011000111111111111111111110100001011111101101011111111100011111111010001111111111001111111111101111111111111111100101111111110101111111101001001011010000010000010000001111111010111111111111111111111111111111110011111010110000111111101001011010000000000000000000000000000000000000000000000000000000000001001010110100000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111111111111111111111111101000010111111011001111111111010111111111010011111110110011101100110101111111111111111011101100111111111111111011000000010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000111111111100011111111110000111111101100111111111010111111111111111111111111111110101111111111000111111110100011000011111111111111111111110000001111111111111111111010111111111011001111111011010111111111000111111110110011100001101011111110101010110000000000000101001011111100001111111010010111111111010111111110101011111111101100101011111111101100111111000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111101100111111111011000001011110111111111111111110101111111110110011111110100101100010100101111111101101111110100101111111111111111111111011000001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010011101111111111111111101011111111101000111111101001011111111101001111111011011111111110111111111111111110101010100101111111111111111111101000000000111111111100111111111010111111111111111110101111111111010111111111000011110100100101001101000000000101000000111111111111111010111111111011001111111110010011111111000011111110110001011111101011111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100101011111111101100111111101000000100111101001111111011011111111110111111111111111111101111010111000101111111110000111111000011111111111111111111111111101100000001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100110011111111110011111111101111111111111111111010111111111101011111111100001111111011010111111110110111111111000101111111111111111111111100000000111111101001011111111101001111111011001111111110101111111111111111110011000000000000000100010100111111101001011111111101011111111010111111111111111111101111111110110011111110100000111111100000111111110001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101101010010111110111111111111111111111111111111111111111111111111111111111111110000011",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010010110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101111111111011111011111111111010000101111101001111111010001111111011010111111110110111111010010011001111111111111011111010001111111111111111111111111111111111110100000001010111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000011111110100101111111110001111111101101111111111011111111111111111111011111111111001011111111000111111110100001111111111111111111111010000101111111111010111111111101001111111010010111111011010111111011010101010000000001001100101111111011111111101100111111101101011111111100001111111011010111111110101111111111101111111011011111110011111111110000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011010100000000000000000100010101010010101111111111111111111111111111111111111111111110100000011",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111101100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111110100111111101010111010000101111111111111111110101111111111010111111111000011111100000001011111110011111111101101011111111111111111111111111111111111111110110100000001001111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010111111110101011111111110100111111110000111111101001011111111101011111111110111110111111111110101111111111000001111111111111111111111011000001101100111111111011111111111111111110111110101010000101010000000001010101000101111111110101111111101011111111111111111010111111111010111111111010001111111110010111111110110011111111010011111111101011111011111100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101101000000000000000000000000000000000000000000010100101011111111111111111111111111111111111011000000111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011111111010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010011111111110100111111101000111100000001011111111011011111111110111111111111111110101111101101010000111110110101111111110001111111111111111111111111111111111111101010110100000000000101011111111111111111111111111111111111111111111111111111111111111111101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000010110111111111101111111111111111111011111111101100111111111101001111111100001111111011001111111110101111110000111111111111111111111110100001010000111111101101011111101101010101010001000000000000000100101111111111000101111110100101111111110000111111101100111111111010111111111111111110111111111110110111111111000011111111000101111111110100111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101000000000000000000000001010101010000010000000000000000000000000100010010111111111111111111111111111100000101111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111101000001111101111111111111111101010111000001101011111111100011111111010001111111111001011111110100011110001101111101011111110110101111111111111111111111111111110101011000000000000000000000000010100111111111111111111111111111111111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111110110101111111110101111111111011111111111111111011011111111011001111111010010111111110010011110001001111111111111111111110110000011011111111101000001011010000000001000000010010101100010111111110101110100101101111111111111111101101111111101000111111101001011111111101001111111010101111111110111111111111111110110011111110110001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101010111011111010101010111011101010110010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011010101000000000000000000000000010101001010101111101111101010101101010000000000000000000000010100111111111111111111110000000011111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111111110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101111111111111111111111111111111110100000111110110101111111101101111111110001001111111111111010111111111011001111111011010111111111000011100010110011111111101011010111111111111111111010101010101101000000000000000000000000000000000000010011111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111110011111111110100111111110100111111101100111111111010111110111111111110101111111011010111110000001111111111111111111111101000010110110101000000000000010100101010111011001111111010010111111111000010100100110011111110101011111111111011111011111111111100111111111100011111111010001111111111010011111110110110101111101111101111111111101100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100010001000100010001000000000000000101010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101010001000000000000000000000000000101010011111111111111111111111111111111111111101110110100000000000000000000010011111111111110100000001111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111000101111111110011111111110101111110100001011111111100111111111010111111111111111110101111111111010110110110100101111110110000001111111111101011010000000100000000000000000000000000000000000000000000000100001111111111111111111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000010101111111011111111101011111111101100111111101000111111111100011111111011001111111110101111111111110000001111111111111111111110110000000000000000010010110001011111111011111111111111111111111111111111001110100101010011111110100101111111110100111111101010111111111011111111111111111011001111111111010111111111000010110110100101111111110011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101000000000000000000000000000001010010111111111111111111111111111111111111111111111111111111111010111101000000000000000001001111111111000001011111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111110000011101111111111111111101011111111000100111111101001011111111101001111111011001111111110101101001110001110111111111111110000111111111011000000000000000000000000000000000000000000000000000000000000000000000001001111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010011111111110011111111101011111111111111111011111111111101011111111100001111111010010111111011000000001111111010101101000000000000000000101101111111101001011111111000011111111010001111111110101111111111000101101111111111110011111111110001111111101000111111111101011111111011011111111110111110111111111110101110101110100011111110100000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000000000000000000000001100000000010011111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000101100000000111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111010010111000011111110110011111111101100010011111111111010111111111011011111111010001111111011000100111010000111111111101111110100101101000000000101010100000000000000000000000000000000000000000000000000000000000000000100001011111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000011111110100101111111110101111111101100111111111010111111111111111010111111111011001111111010000000010101000000000000010100101010000101111111111111111011111111111010111111111101001111111010010111111111000101111110101011111111111111111111111111101101111111101101011111111100001111111010001111111111001111111110110111111111111111101011111111110100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000000000000001010100101111101100010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101000000000000010000000100111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100010100110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111101111111111111111111111111111111100010110110111111110100101111111110000001111101100111111111011111111111111111111111111111111000001111100010011111111000011000011100000000101011111110000000000000000000000000000000000000000000000000000000001010000000000000101001111111111111111111111111111111110110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000101111111101111111111110101111111110001111111101001011111101101011111111010111110111010101100000000000000010101010010111111111110100000111111110100111111111010111111111110111110111111111011001111111111000011111111000011111110110101111111101011111111111011111111111111111010111111111011001111111010010111111111000011111110110011111111101011111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010000000000000101010111111111111011000101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101000000000000000000011111111111",
"0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111110111111111111111111111111111111111000010111111111111111111111111111100001011111101000111111101001011111111101011111111110101110110101101000101111111110110100000100000001001111101100000000000000000000000000000000000000000000000000000000000000010100000000000000000100101111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111110001010111111110101111111111111111111011111111101100111111111001011111101100010101000100000000000000000010101111111111111111111111110001011111110100111111101001011111111101011111111010111111111111111110100101111111101111111110110101111111100100111111110100111111111100111111111110111110111111111110101111111111000011111110100101111110100101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000100101011111111111011010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000010111111111111",
"0000101001010110010101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111010101111111111111111111111111111111000010111111110110011111111101111000100111111101011111111101010111111111101001111111100001110110011000101111110101110110101010000010011111011000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100101111111111111111111111111111111111111010010111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111010000011111110100011111111110101111111101011111111111011101101001101010000000000000000010101001100010011111111111111111111111111101000010111111011111111101101111111111101011111111100001111111010001110100011001111111111111111111111111111101011111111101000111111101001011111111101001111111011011111111110111111101011111110101111111111110101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111111111111111111111111111111111111111111111111111111111111111110110100000000000000111111111111111011010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000001001111111111111",
"0101010101100101010101010101011101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101101111111111111111111111111111111101100010111111111010011111110100101000101110101111111101011111111111111111110111111111111001111010010000011111111000101010011101101111010100000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000100111111111111111111111111111111111011010111111111111111111111111111111111111111111111111111111110110111111111111111111010111111111111111111111111111111111111111111111111111110110000111110110011111110110101111111110000111011010100010000000000000000000101001110111111111110010111111111111111111111111111101100000101111111101011111111111111111011111111111010111111111011010111000100010111111111000011111110110011111111101111111111111111111010111111111101011111111010010111111011010011101101010111111111101011111111111111101000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111101100000000000000010111111111111010110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111",
"1111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110011111111111111111111111111111111101000001111111111101111111110110000000101110100111111101000111111101100101111111010111111111011001111010011111111001011111111111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010100111111111111111111111111111110010111111111111111111111111111111111111111111111111111111111010111111111111111111011011111111111111111111111111111111111111111111111111111111100001111111111111111101011101010110000010000000000000000000000010101101001001111111011001111000011111111111111111111111111111100000101111111110000111111101100111111111010111111111110111111111110100010101111111111010111111110100011111111110101111111101101111111111011111111111111111010111111111111010111101000000011111111000101111110110101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111011010000000000000101011111111111111100001010101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111001111111111111111111111111111111110100001011111010111111110101111111100000111111011111111101010111111101000111111111100011111111100001111010010101111111111111111101100000000000000000000000000000000000000010101010011001101010101000001000000000000000000000000000000000100000100000000010000010011111111010011111111111111000011111111111111111111111111111111111111111111111111111111000111111111111111111101011111111111111111111111111111111111111111111111111111111111000100111110100101010100000000000000000000000000000000000000000100010000010010111100001111000101111111111111111111111111111111000101111111101011111111101000111111101001011111111101001111111010000111111110111111111111111110101011111111110101111111110000111111101001011111111011011111111110111111111111111100001111111110110011111110100100111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110110000000000010101010011111111111111101010110011010101000000010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111011011111111111111111111111111111111111000001011011010111111111000011111000000011111111101011111111111111111111111111111010111111111100001110001010010111111111111011000000000000000000000000000000000101010010101111111111111111111111111010101011010101000000000000000000000000000100000001001011000000010010000101111111111111000101111111111111111111111111111111111111111111111111111111000111111111111111111100011111111111111111111111111111111111111111111111111111111111110000010100000000000000000000010101000000010101000000000000000000000000000001000000010011000101111111111111111111111111111110100000110011111111111011111111111111111010111111111101001111111010000011111110010111111110110111111111101111111111111111111011111111101100111111111001001111111100001111111011010100001110101111111111111111111011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111101100000000000101111100001111111111111111111111111111111111111110110100000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101010101110111010111010111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111111111111111111111111111111100000001011111111111111110101011101000000011111111100101111111110100111111111100111111111011101100111101001011001111111110110000000000000000000000000000000101010011111111111111101010101111111111111111111111111111111111010000000000000000000000010000000011111101000000000001111111111111000100111111111111111111111111111111111111111111111111111111000111111111111111111100001111111111111111111111111111111111111111111111111010110100000000000000000000000001000101001010110001001011010001001011010000000000000000000000000000000000101111111111111111111111111110110000000101111111110100111111101100111111111011111111111111111011000011111011001111111111000011111110100101111111110101111111101011111111111111111110111111111011001111111010010100001111000111111110100011111111110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111000000000000000100110101111111111111111111111111111111111111111111111010110000000101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101101010101010101010101001011001011001100110010110011001010111010101010101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011101101111111111111111111111111111111101100100001001111111110101111111111110001001111111111101011111111101100111111101001011111111100010101101100001100111110101101000000000000010000000000000001010011111111111111101101000000001111111111111111111111111111111111101011000000000000000000000000000000111110101001010001001111111110100000111111111111111111111111111111111111111111111111111111000011111111111111111100010111111111111111111111111111111111111111111010110000000000000000000000000000000100000001000000000000000000000000010101000000010101010000000000000000000001010011101111111111111111111111101000000011111111110100111111101000111111101001011111111101011111000010111111111111111110111111111110110011111110110101111111110000111111101100111111111010111111111111111110111010010111010111111111000011111110100101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111111111111111111111111111111111111111101000000000000000000000000101111111111111111111111111111111111111111111111111111111010000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111110111011101010101010101010101010101011101010101011001010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101011111111111111111111111111111111110010100000001111111010010111111111000000111111110011111111111011111011111111111010111111111100000011110000000010101100000000000000000000000000000001010010111111111111101101000000010011101111111111111111111111110100111111111111101101000000000000000000000000010111111110111010010011111111110001001111111111111111111111111111111111111111111111111110100101111111111111111010010111111111111111111111111111101110101101000000000000000000000000000000000000000000000100000000000000000000000000000000000000000101000000000100000000000000000001010100111111111111111111111010010111101111111111111111101011111111111100111111101101001111000000001111111111010111111110101111111111111111101011111111101101111111101001011111111001011111111011001111111010000111111111111111101111111111110011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111111111111111111111110100000000000000000000000000001111111111111111111111111111111111111111111111111111111111011000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101101111111111111111111111111111011001110000001111111111110101111111111000101111110100011111110110101111111101101111111111011111111000010100000001111000000000000000000000000000000000100101111111111101101000000010010111111111111111111111111111111101100000010111111111110101100000000000000000000000101011111111111000100111111101000010111111111111111111111111111111111111111111111111110100101111111111111111010010111111111111111111010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000010011111111111111111010000010100101111111110101111111111011111111111111111010111111000101001111111010010111111111000111111110110011111111101011111111111111111111111111111011011111111100001111111010000111111111000111111110110011111111101011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000010011101111111111111111111111111111111110111011101111111111111111101101000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111101011100000101111010101111111110111111000011111111101011111111110101111111110100111111101000111111000101000001001010000000000000000000000000000001001111111111101101000000000100101111111111111111111111111111111111111100000001010111111111111110110000000000000000000000010110111111101000011111111100010011111111111111111111111111111111111111111111111110100001111111111111111111000011111111111010110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010100001010011111111111110100100110011111111110100111111110000111111101100111111111010010111111111111110111111111110110111111110100011111110100101111111110100111111111010111111111111111110111111111011000111111111010011111111000011111110100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111110000000000000000000001000001001010101111111111111110111010110101010101010101010101010100101011111110101100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111110101111100000101111100001111111010010111000010110111111111101111101111111111101011111111101100111111010000000001010000000000000000000000000001010011111111111011000000000000010111111111111111111111111111111111111111111100000000000101011111111111111111010000000000000000000101001111111100010111111010000101111111111111111111111111111111111111111111111111100000111111111111111111000000101101001000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100101011000101001111111110100001011111111111101011111111101101111111101101011111111000010011111011001111111110101111111111111110111111111111110011111111110100111111101001011111111101011111111011011111000100111110101111111110110011111110100101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000100110010111111101010110101010101010011001100101010110101010101010101011111111011110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111110100101111010000101111111011111111011010111000011000111111110100011111111110011111111101011111111111100010100000000001100000000000000000000000100111111111111110100000000000000010111111111111111111111111111111111111111101000000000000000010011111111111111101100000000000000000000010111101000000011111111000000111111111111111111111111111111111111111111111111110000111111111111111111000000000000000000000100111010000000000000000000000000000000000000000000000000000000000000000001000001000101000100000000000000000000000000000000000000000000000000000000010011111101010100111111101000001110110011111111101011111111111111111010111111111010010111111100001111111010010111111111010111111110101011111111111111111011111111101010111111101101011111111100001110100001010111111110110111111111101111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111101100000000000000000000000100000001011110101101010101010010111011111111111111111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101010100110011001100110010101010101111101010111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111011000001011010000100111111111110111111111010010110101111111110110011111110100101111111110001111111101001001000000001001100000000000000000001001111111111111101000000000000000000010011111111111111111111111111111111111011000000000000000000000000111111111111111110110000000000000000000011111100000101111111100001011111111111111111111111111111111111111111111111110001001111111111111110101000000000000001011110110000000000000000000000000000000000000000000000000000000101010100101010111110111010111011111010101100110101010000000000000000000000000000010000000001001111101100010111101000010110100101111111110001111111101100111111111010111010010011111110111111111011001111111111010011111111000011111110100101111111101011111111111011111011111111111010101110100000001111111110010011111111000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111110110000000000000000000000000000010010101101010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010010101011001010101010101010111010101011101011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111011010101011010000000011111111100001111111010010011111110101111101111111111101111111111101101111111101001010000010000000000000000000000010101111111111110110000000000000000000000000000111111111111111111111111111010110000000000000000000000000000010111111111111111101011000000000000000001001010000101001111101000001111111111111111111111111111111111111111111111111000001111111111111111111001010000010011101101000000000000000000000000000000000000000000010101010011111011111111111111111111111111111110101011001101001010111111101011010000000000000000010000000000000100111111000001010000000011101111111111110010111111110000111111101001011111000101011111111010111111111111111111101111111110110111111110110101111111110000111111101000111111111100111111111110100000111111111110101111111111010011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000010011111111111111111010000000000000000000000000000001010011010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111101000111111111010000101111111111011001111111100010111111111010111111110110011111111101111111111111111110001000001001000000000000000000100101111111111111010000000000000000101000000000000010111111110111111111111010000000000000000000000000000000000010011111111111111111110110000000000000000010011010011010011101000000100111111111111111111111111111111111111111111111010010111111111111111110101001001001111101010101010100000000000000000000000000000010011101111111111111111111111111111111111111111101100000000000000000101010101111111111010110100000000000000000000000000010010100001000001000101111111101011111111111111111011111111101100111111000001011111111100001111111011010111111110101111111111111111101111111111101011111111101100111111101001011111111100000001111011001111111110101111101111111110110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000101111111111111101100000000000000000000000000000001010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111100000111111101100000011111010111110111111101001001111111111010111111110100011111110100101111111110100110101000001010000000000000001010011111111111111111100000000000000000000000000000001001111111101010111111011000000000000000000000000000000000000000101111111111111111111111011001011010000000001000000110111111010110101010100111111111111111111111111111111111111111010000011111111111011000101000011111111111111111111000000000000000000000001001010111111111111111111111111111111111111111111111111111100000000000000000000000000010100111111111111101011000000000000000000000000000110101100000000111110100101111111110101111111101010111111111010001110111111111010101111111011001111111110000111111110100011111111110011111111111011111011111111111010111111111101000000111010001111111011010011111110110011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000100000000000000000101111111111110100000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111110100011111111101000000011101101011111111011010001011110111111111111111110101111111111110011111111110001010000000000000000000000000010111111111111111111101000000000000000000000000000000001001111101101010111101100000000000000000000000000000000000000000001011111111111111111111111111111101001001101010001001011111111111011101101010000001111111111111111111111111111111110100000111111111011001010111111111111111011101100000000000000000001001110111111111111111111111111111111111111111111111111111111111111101011000000000000000000000000010011111111111111101011000000000000000000000100111011000000011110110011111111110101111111110000111111101001001111111010111111111111111110111111111110101111111111010011111110100101111111110100111111101101111111111011111111110001011010101111111111010111111111000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000111111111010000000000000000000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111011011111111111111100000101111100111111111101000100111010010111111111010111111110101111111111111111101010000000000000000000000001001111111111111111111110110000000000000000000000000000000100111111101010111111110000000000000000000000000000000000000000000001001111111111111111111111111111111100010110111100001111111111111111111111101101001111111111111111111111111111111111110100111111111011111111111111111110110000000101010000000000010011111111111111111111111010111111111111111111111111111111111111111111111111110000000000000000000000000001001111111111111110110100000000000000000000010111101000010111111111111111101111111111101101111111101001011111111000011111111100001111111111001111111111101111111111111111101011111111110101111111110000111111101101001111101000011111111110111111101111111110101011111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001010000001001111101000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111100111111110101111110000101111111111011111110110000111011011111111111010111111111010011111110110101111100000000000000000000000101111111111111111111111010000000000000000000000000000000000011111110111111111111000000010000000000000000000000000000000000000000010111111111111111111111111111101001010111111011000011111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111110110101001110100001001110111111111111111111111011000101011111111111111111111111111111111111111111111111111000000000000000000000000000000100111111111111111011000000000000000000000101111010000101111110100011111111110011111111111111111111001111111010111111111011001111111010010111111111010111111110110111111111111111111111111111111010111111111101011111101000001111111010010111111011010111111110101111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001010000000000001110100000000000000100000000010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111110011111111111111111111101001111111110001111111000000111111111101011111110001011111111111111110101111111110110011111110100100101000000000000001000000001111111111111111111111101000000000000000000000000000000000000011111111111111111100010010110000000000000000000000000001000000000000010011111111111111111111111111110101101111111110110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111000100111111111111111111111111101100000000111111111111111111111111111111111111111111111111101000000000000000000000000100000001001111111111111111101100000000000000000001011111000100111110110011111110100101111111110000111111001100111111111111111011111111111110111111111111010111111111000011111110100101111111110101111111111011111111111111111100001111111011001111111110010111111111000011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000001000101000000010010000000000000010000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111110110111111111111111111111110011111111111011111011000000111111101101011111110000001111111011001111111110101111111111111110100000000000000000000000000100111111111111111111111011000000000000000000000000000000000000000100111011000100110000010011000000000000000000010100000010101101010000000101111111111111111111111110110011111111111111101100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111110100000000101111111111111111111111111111111111111111111111111100000000000000000000000010100000000000100111111111111111011000000000000000000000011100001001111101111111111101011111111110100111011010001011111111001011111111011011111111110111111111111111110101111111111110011111110110001111111110000111111101100111100010110111111111111111110111111111111010011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000010011000000000100000000000001010000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111110101111111111111111111111010011110101111111101100000011111111111011111110110001011111111011010111111110010011111111010011101010100000000000000000010011111111111111111111101100000000000000000000000000010000000000000001010000000000000000000000000000000100110000010101010101010111101000000101111111111111111111111111010111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000010111111111111111111111111111111111111111111111111110100000000000000000000000000001010000000000001111111111111111111100000000000000000000101000000111111110110111111111101111111111111101001011111111101101011111111100011111111100001111111111001111111111101111111111111111101011111111101101111111101001011010010000011111111011001111111110101111111111111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100110000000000000000000000000101000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111011001111111111111111111111001110110101111111110000000101101100111111111011000100111111111110111111111010101111111111010011111111000000000000000001001111111111111111111111110000000000000000000000000100110000000000000001000000000000000000000000000000000010100000000000111110000011101011000000111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111110101100000000010111111111111111111111111111111111111111111111111101000000000000000000000000000000000000000000000100111111111111111110110000000000000000010100000011111110100011111110110101111111101001011111101011111111111111111010111111111011001111111011010011111111000011111110110011111111101011111111111111111011111010000101011111111100001111111010010111111111010011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000101000000000000000000000000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111011001111111111111111111100001111101111111111101101000101101000111111101000000101111101001111111111011111111111111111111111111010010000000001000000111111111111111111111110100000000000000000000000000100110000000000000000000000000000000000000000000000000000010011110000001110101010010110100000111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111011000000000000000101111111111111111111111111111111111111111110110000000000000000000000000000000000000001000000000001001111111111111111111100000000000000000000000011111110101011111110110101111110100000111111101000111111111100111111111010111111111111111110101111111110110011111110100101111111100101111111101100111111111100000011111111111110111111111111010111111110000111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100111111111111111111111100010011111111110011111111000100111111111111111101000101111101011111111010010111111011010111111110110101010000000000000101111111111111111111111110100000000000000000000000010100000000000000000000000000000000000000000000000001000000000111110000000000111111000010100000111111111111111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000010011111111111111111110100000000000000000000001001111111111101111111111111111110000111111101100111111101001011111111101001111111011001111111110101111111111111111101111111111101101111111110000111111101000000011111101001111111010101111111110111111101111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001001100000000010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111100111111111111111111101001000011111110100101111110100001111111101011111111000101111111111111111010111111111111010111111111000000110000000000000011111111111111111111111111000000000000000000000000010000000000000000000000000001000000000000000001000001010010010010000100110000101010101011000001111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000101010100101110101111111111111111101100000000000000000000000000000000000000000000000000000000000000111111111111111111101100000000000000000000000111111111000011111110110100100000101011111111111111111011111111111101011111111010001111111010010111111111010111111111101011111111101111111011111111111100000101101100011111111100001111111011010111111110101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100101000010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111101100111111111111111111110101111111111111101011111110100001111111110000111111000001011111111010111111111110111110111111111110100100110000000000010011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000101000000101010111100000111101100110000111110000101111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000100010111111111111111110000000000000000000000000000000000000000000000000000000000000001001111111111111111111111000000000000000000000100110100000111111110100100100101100100111111101100111111111011111111111111111110111111111111001111111111000111111110100011111110110100111111101011111110100101111110111111111011011111111010010111111110000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010100001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111101101111111111111111110100111111110101011111111111111110000111111111101111111000001011111111100001111111011001111111111001111110100100000000000010111111111111111111111111100000000000000000000000000000000000000000000000000000000000001000000010101000100100000111011001010010111110000101100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000010011111111111111111111101000000000000000000000000101001111111111101111000101110101111111110000111111101001011111111101011111111010111111111111111111101111111110110011111111110101111111110000111111100001011111111010111111111110111111111111111010101011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001001100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111110011111111111111111111010111111111000011111110100011110000101101111111111011000011111111111010111111111010001111111010010110100011000000000000010111111111111111111111111000000000000000000000000000000101000000000000000000000000000000000000000000010011110100111111101100010010101110110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000000000000000000101111111111111000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111011000000000000000000000111111110110011111111000101111111111111111011111111101100111111111101001111111100001111111110010111111110101111111111101111101011111111101101111111110001011111111000011111111100001111111111001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111110110011111111111111111011001111111110101111111110110101110001000101111111101000000011111100111111111010111111111111111110101110010100000000010100001111111111111111111111101000000000000000000000000001001010100000000000000000000000000000000000000000001111111011111111101001001010010111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000100111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110110000000000000000010111111111000011111111000101111111110101111111101011111111111111111010111111111010101111111011010111111111000011111110110011111111101011111111111011110001011111111010111111111011001111111010010111111011010010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111110110111111111111111111101011110101111111111101111111111101000001011111111101000010011101001011111111101011111111011001111111010010100000000010101001111111111111111111111110000000000000000000000000000001110100101000000000000000000000000000000000101111111111111111111101001111010010011010000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000000000000000000000000000000010010101100000000000000000000000000000000000001000000000000000000000000000000000001011111111111111111111111111100000000000000011111111111101111111010000011111111110101111111110000111111101101011111111010111111111111111110101111111110110111111110100011111110100100111111110100101001011100111111111011111110111111111011001111111111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111001111111111111111111100111010010111111111010011111110110001011111111011111010000011111010111111111101011111111100001111111100000000000000001101011111111111111111111110110000000000000000000000000000001101001111000000000000000000000000010101010111111111111111111111101100101010111010000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011000000000000010011010011111110110010010111111111101011111111101010111111101000111111111001011111111100001111111110101111111111111111101111111111101011111111110100111000010001011111111101001111111011011111111110101110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111001111111011001111111111111111101000111110101111111111010011111110100000001110110101111111000100111111111011111111111111111110101111111100000000000000001001011111111111111111111011000000000000000000000000000001001000001110101011000000000001000000010111111111111111111111111111111110100001111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000010111111111111111111111111110100000000000000100010111111111000000001110110011111111101011111111111111111111111111111010111111111011001111111010010111111111010011111110110111111111101111111011111100000010111111111101011111111100001111111010010111111111010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111110111011101110101010101010101010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111011111111010111111111111111111111001001111111111111111111111111111101100001111110101111010000000111111101001011111111101011111111010101000000000000001001000111111111111111111111111000000000000000000000000000001111101001100001110100101000100101100001111111111111111111111111110111111110001110000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000001000000000000000000000000000000000111111111111111111111111111101000000000000000001111111110110001001110100101111111100100111111110100111111101010111111111110111110111111111110101111111111010111111111000101111111110101111111101000010111111011111110111111111010111111111011001111111010000101001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110111010101010101010101010101010101010101010101010101010111010111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001111111111111111111111111111111111111111111010111111111010111111111111111111101000001111111011010111111110110111111010010111111111111111000101111111111100111111111101011111111100000000000000000000110000111111111111111111111110100000000000000000000000000100110011101000001010101010100101111101001111111111111111111111111011010010110010100000000000000001011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010001001000010000000000000000000000010111111111111111111111111111111100000000000000001110101111101101011111111111111111101011111111110100111111101001011111101101001111111010101111111111111111101111111111101111111110110101111111110000000111101000111111111100111111111110111110111111111110111010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101101010101010100110100110011011010111010101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110101011101011111111111111111111111111111111111111111111111111111111111111010011111111111111111111111111111111111111111011011111111010111111111111111111101001011111111111001111111111010011111010000011111110110100010111101011111111111111111010111111111011000000000000000001010001111111111111111111111110100000000000000000000000000011000101101010101100001110100100100011111111111110111011010101010000000000000001000000000000000000010000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000010101000100110000001011010000000000000000000000000011111111111111111111111111111010000000000000000100010111111000000011111110101011111111111111111011111111101010111111111101011111111100001111111010010111111110110111111111101111111111111111101100000011101000111111101101001111111100001111111011010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110101010101010101010101010111110101010111110111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111101111111101101111111111111111111110101111110111111111111111110101111111111000011111111110000010111110001111111111100111111111010111110100000000000010001000101111111111111111111111111100000000000000000000000010010000011000101101001001101001111000000110101010100000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010101001100001100000100110000000000000000000111111111111111111111111111111111000000000100000000001111101000010111111110100011111111110101111111101011111111111011111110111111111010101111111011001111111110010011111111000011111111110011111010000101111111111111111010111111111101011111111100001111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010101010110010110100101010110010110010111011101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111101101111111111111111111110100111010001111111011001111111110101111000011111111101010010111101101111111101001011111111100011111000000000000000000000100111111111111111111111111110000000000000000000000010000011111000100101010110000010101000000000000000000000000000000000000000000000000000000000000010001001010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000001000100000000000000000000000000000000000000000000000100000000000101101000010000000001000101101000000000000000000011111111111111111111111111111110100000000000000000001111101000111111111110101011111110110101111111110000111111101001011111111100111111111110111111101111111111101111111110110011111110100101111110000001111111101100111111111011111111111111111110101111111011010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101100101100110011010101001100101010101010111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111110011111111111111111111110001111011011111111011010111111111010110110010110011111011000011111111111111111011111111111100111011000000000000000000000101111111111111111111111111110000000000000100010101010001001010110011000101010000000000000000000000000000000000000000000000000000000000010101001011111111111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000010000000000000000010000010100000000000000000000000000000000000001000000000000000000000001010100000001000001101011001100000000000000000101111111111111111111111111111111101000000000010001001011000100111110110111111111101111111111111111101011111111101100111111101101011111111100001111111111001111111111101111101111111111101111111111000001111111110000111111101101011111111101001111111010111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110111111101010101010110101010011001100101011001010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110101111111111111111111111110000111111111111111110111111111111010111100000100011111110000101111111110100111111111010111111111010000100000000000000000000111111111111111111111111110000000000010010000101101001010000010100000000000000000000000000000000000000000000000000010101010100101100111111111011111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000000000000001010100000000010100010001000000000000000000000000000000000001010001001100000000000101000100111100010110110000000000000000111111111111111111111111111111101100000000010001011111000001111111000111111110100011111111110011111111111011111111111111111010111111111011001111111010001111111011010011111110110011111111101010100000111111111010111111111100111111111100001111111100010111111011010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111110101110101011001100110101010101001100110010101010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111110110111111111111111111111110001011111111011001111111110111111111111110000101111111111000011111111110001111111101001011111111000010000000000000000000100111111111111111111111111110000000000010111000101010001010000000000000000000000000000000000000000000100010100101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100010000000000000000000000000000000101101000001111000000000000000000000000000000000101111100010011010000000000000001010100001110110000000000000000111111111111111111111111111111111011000000010100001110100100111110101111111110110011111110100101111111110001111111101100111111111011111111111111111110111111111111010111111111000011111110100100100001010101111111111011111111111011111011111111111011001111111010010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111010101010101100110101010101010101010010110010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111110101111111111111111111111100101011111111010001111111010010111111010000001011110101011010111101111111111111111101101111111101000000000000000000001000000111111111111111111111111101000000001010100000000000000000001000000000000000000000000000000000101010011111111101011111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010100000000000000000100000000000001010001001111000100101100000100010101000000010010101100010111100000100001001100010111110100110001000000000001011111111111111111111111111111111110100000000000010111100001001111111110101111111111111111101011111111110101111111101000111111101001011111111011001111111010111111111111111111101111111111110011110000000100111111110000111111101100111111111010111111111111111110111110100101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101010101010101001010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111011001111111111111111111110110101111111111011111111111111001111111010000000011110100011010110110101111111101011111111111011101001000000000000000000000001001111111111111111111111111100000000000000010100000101000100000000000000000000000001010100101111101111111111110011111111101100111111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010000000000000000000000000000000000010100110101111100001010101011000101001100010011001110100000101000010011010110110000101011000000000001011111111111111111111111111111111110100000000000010011100000010111111111010111111110110011111111101111111111111111111010111111111100111111111100001111111010010111111111010111111110101111111111110000001011111111101100111111101001011111111000001111111100001111111010000100101100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111011111111111111111111110100011111101011111111010111111111111111010000011001110110011010111110101111111110001111111101100110000000000000000000000000000001111111111111111111111111110000000000001001101000000000000000000000000010000010010101111111111111111111111111011111111111010111111111010111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010100010000000000000000000000000001001101010100001110100000101010101100010111110000101100111100000010101101010000111010000000000001011111111111111111111111111111111111110000000000000010110100101111111111010111111111000011111110100101111111110101111111111010111111111111111010111111111011001111111011000111111111000011111110100000011111101011111111111111111011111111111010111111111100001111111010000000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111011011111111111111111111110100111111101011111111100001111111110001111000011010110111110010011101111111111101101111111101001010000000000000000000000000100010011111111111111111111111111000001000001000000000000000000000001010100101111010111111110101011111111110111111111101011111111111011111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101000000000000000000000000000100010111110100110100111100010010101011110000111010010011000001000001011111010011010000000001011111111111111111111111111111111111110000000000000000000111111110111111111111111111101111111110110011111111110001111111101000111111101100111111111010111111111111111110111111111110110111111110100000001111100100111111110000111111111100111111111011111110111111111011010001011111010010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100111111111111111111111110100011111011111111111010111111111011010111000101000010111010000011111111101011111111101111111010100000000000000000010001000000110011111111111111111111111111100000000100000000000000000101010010101111111110101111111110110111111110110011111111101011111111101010111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101011010100000000000000000010110000101011001010010111110101101010101111010111100001001100111010000011101100000001011111111111111111111111111111111111100000000000000000010011111010001111111111010111111110101111111111111111101011111111101100111111101001011111111101001111111011010111111110101111111111111111101000010111110011111111101100111111101001011111111101001111111011011111111100010110101111101011010000000000000000000000000000000000010000000000000000000000000000000000000000001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111101101111111111111111111111111000000111111111010111111111110111110111111000100101100111100000011111110100101111111110001111111000000000000000000000100110101111111111111111111111111111111101000000101000000010000101010111111111110111111111111111111111111111111111011111111101111111111101011111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101101010100000000000000000000111010000110101101101011111110101111111111110001011011010101010011110000000001011111111111111111111111111111111111110000000000000000010111111011001111111011010111111111000011111110110011111111101011111111111111111110111111111011011111111010001111111010010011111111000011111100000011111111101111111011111111111010111111101101011111111100001111111100010111111111001111101011000000000000000000000000000000000000000000000000000000000000000101010000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111101011111111111111111111111111000000111111111001011111111101001111111111000101111101001100010111111111101011111111110101111111000000000001000001010001011101111111111111111111111111111111101100000000010101001011111011011111111010101111111111001111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111110110100010000000000000001010010010111110000111111111111111111111111101000001110000011101101010000000001011111111111111111111111111111111111110000000000000000010010111111111111111110111111111110110011111110100101111111110001111111110100111111111010111111111111111110111111111111001111111110110011111010000011111111110101111111101010111111111011111010111111111011011111111010000101111010000111111111000100101100000000000000000000000000000000000000000001010101001111111100010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111101011111111111111111111111111010011111111101010111111111011001111111010000101101100000000010110101111111111101111111011111100000100000000000101111100001111111111111111111111111010101010101101010011101111111111111010111111111110101111111110110111111110110111111111101111111111111110111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111110111110110011010101010000000000000011101100101011111111111111111111111111101100000010110011101000000000000001011111111111111111111111111111111111110000000000000000001100001111111011001111111110101111111111111111101111111111110011111111110000111111101001011111111101001111111010101111111110111110101111111010000011111111100101111111110001111111101000111111111100111111111010111110100100111110101111111111010011111111000100101101000001010100000001001011000100111011111111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111110111111111111111111111111110010111101101111111111110111110111111111111000101101000010001001111000011111110110101111111110100010010000000000011111111010111101011111111110101101101010101001011111010111111111010111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111110101111110001001011000000000001010001011111111111111111111111111111111011000101101100001100000000000001011111111111111111111111111111111111110000000000000000011011011111111010001111111011000111111111010111111111101011111111111111111011111111111100111111111101011111111010001111111111010111111110101010000011101111111111101111101101111111101101011111111001011111111100001111110001001111111110101111101111111111101011111111110100111110100000101110100001011111111101011111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110110111111111111111111111111010001111101000111111101101011111111011011110100100110000111101001110101111111111100011111111110000001100000101000011111111101111101111111111101010111010101101111111101010111111111010111111111010101111111110101111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111110101010100000101000000000001011111111111111111111111111111111110101010101000001111000000000000111111111111111111111111111111111111100000000000000000001111111111111110111111111111001111111111010011111110100101111111110101111111101011111111111111111010111111111011001111111010010111111111000011000100100011111111101011111111111011111011111111111010111111111101011111111000010111111010010111111111010111111110101011111111111111100001011110110000111111101000011111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111001111111111111111111111111100010111111010111111111101011111111100001110100000000101111100001111111111101111111111111111110000001100000100010111111111111111111111111111111111111111111111111111111011111111111010111111111111011111111111001111111111101111111111111111111110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011101100010010110000000001010111111111111111111111111111111111111100001010101010000000000000111111111111111111111111111111111110100000000000000001011111111100011111111010101111111111111111101111111111110011111111100101111111110000111111101001011111111010111111111111111111111111111110101111000101010011111110100101111111110001111111101100111111111011111110111111111100001111111111010111111111000011111110100101111110110101101000010011110000111111111010111111101000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111110111111111111111111111111111010010101111111111011111111111111111010111111100000000001111010010011111111000011111110110011110000010000000100001111111110110011111110110011111111101101111111111011111111111111111111111111111111111111111111111111111110111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010101001101010000000100111111111111111111111111111111001000011110100000000000000011111111111111111111111111111111111111000000000000000001011111111101001111111100010111111111010111111110110111111111111111111011111111101010111111101100111111111001001111111100001111111111001111111111000001101111111111101011111111110101111111101000111111101001011111111101011110010010101111111111111110101111111110110011111110100101101000000000101000101000111111111010111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001111111111111111111111111111111111111111111111111111111111111111111111111111001111111111011111111111111111111111111010000100111111101000111111101100111111111011000100110000111010001111111110110011111110100101110000000000010000001110101110101111111111101011111111101101111111101101111111111111111111111010111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111010111010100101010001000000010011111111111111111111111100001110101011000000000000000011111111111111111111111111111111111010000000000000000000111011111110111111111010111111111011010111111111000011111110100011111111101101111111111111111011111111111010111111111011001111111010010111111111000100111110110011111111101111111011111111101011111111111101011111111100001110100000001111111011010111111110101111101111111111101011111010000001111001010001011111101001001111000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111011011111111010111111111111111111111111111100010011111111101101111111111001011111111100000101101001001011001110101111111111111111101110100001010000010101001100001111111111111111111111111111111111111111111111111111111111111111111010111111111011111111111010101111111110101111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111110110011010101101100000000001111111111111110101100001110100000110000000000010011111111111111111111111111111111111010000000000000000001101101011111111010111111111111111111111111111110101111111110110011111110100101111111110000111111111100111111111011111110111111111110111111111111000000111111000011111110100101111111110101111111101011111111111111111011111111110000001111111010010111111110000011111110100011111111110100000100111100001011111111111100111110100000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111111111010111111111010111111111111111111111111111100011111111011111111111111111011111111111010000101110000001010001110010111111110110011111111000000110000000001010011010111111110110011111111101011111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111101111111111101111101101010101010000000100101111111010010110110100100001000000000000010111111111111111111111111111111111111010000000000000000101101101011111111000011111111100001111111010101111111111101111111111111111101011111111101100111111101001011111101100011111111011011111111110111111110001011111101111111111110011111111110001111111101000111111111100111111111010101001011111111110111111111110110111111111000011111110100001000000110000001111101010111111111011111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111101111111111111111111111111111000001111110101111111101100111111111010111110100101101001011011010111001111111111010011111111000101000000000000111111101111111111101011111111110011111111111111111111111010111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111101011111111111111101100101101010000000000000010111101001110110000101100000000000000001111111111111111111111111111111111111100000000000100000101111011111111111010111111111011001111111110010111111111010011111110110011111111101111111011111111111011111111111101011111111100001111111010010111110000010111111110101111111111111111101111111111101100111111101001011111101100011010001011001111111110101111111111111111101111111111110010100001010000010111110000111111101101011010000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111111111111111101111111101101111111111111111111111111101001011111110101111111110100111111101001011111100001010100111010010111111111111110101111111110000100100000001000111111111111111111111111111111111111111111111111111111101111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111010010010100000000000010010110100110101101100000000000001001111111111111111111111111111111111101000000000010000000000111111101010111111111011111111111111111110101111111111010111111110100011111110110100111111101101111111111011111111111111111110111111111011001111101000000111111110100011111110110011111111101011111111111111111011111111111101001111010100001111111010010111111111010011111110110111111111110000001011010011101100111111101001011110100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011101111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111101010111111101011111111111111111111111111101000010011111111111111111011111111111100111110100000010001011010010011111111010111111110101010000101000001011000001111111110101111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111101100111111111111111010101110110000000000000001000001011011010000000000000001011111111111111111111111111111111111110000000000000000000100111111101001011111111100011111111011001111111110111111111111111110101111111110110101111111110001111111101000111111111100101111111011111111111111101000001111111110110011111110110101111110110100111111101100111111111010111111010111000010111111111011001111111111000111111111000011111110100000001111000101111111111111111111111111101000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101101001010101010111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111110011111111111111111111111111101000000011111111110101111111101011111111111110100100101000111011000011111010010111111111000000000100000000111100101111111110110111111110110011111111101011111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111011111110111111111111111111110010110000000000000000010100000000000000000101111111111111111111111111111111111110100000000000000000001111111111111011111111111101011111111100001111111011010111111111010111111110101111111111111111101011111111101100111111101101011111111100001111111011000000001110101111111111111111101111111111110101111111110000111111101001011110100000000101111010111111111111111110111111111110110011101110100000000111100001111111101000111111111100111110000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010101101001100110010101111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111110111111111111111111111111111110000010011111111110100111111110000111111101100000011110001011110100101111111111111111110110000000000000001111111111111111111111111111111111111111111101111111111101111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111001111111111111110101111111011000000000000000001000000000000010111111111111111111111111111111111111111000000000001000000011111101101111111111011111111111111111010111111111011010111111111000111111110100011111111110011111111101011111111111111111010111111111011001111111010010000001110010011111110110011111110101111111111111111111111111111101010111111101001001000111100001111111011010111111111001111111111101111111010000101110001111111110100111111101001011111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111010101010101100101111111111111111111111111111111111111010101110110101010100110111101111111111111111111111101011101010101011111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111111111111111111111110100100010111101111101011111111101101111111101000000011110001001111110000001111111110101111111100000000000101111111111110101111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111110011111111111111111010110000000000000000000000000001011111111111111111111111111111111111111010000000000001000001011111110000111111101101011111111101011111111010111111111111111110101111111110110011111110100101111111110100111111101101011111111010111111111111111110111100010110110111111111000011111110100101111111110101111111101011111111111111111100011100111011011111111010001111111110000111111110110011111111000101101001011011111111111111111010111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111110111010101101010100110010101011111111111111111111111111111010101011010101010010101110111111111111111111111111111010101011001100110010101111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111110100100001110110011111111101011111111111111111011000111110001011111110000001111111110010111111100000000000011111111111111001111111110101111111111111111111111111011111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111110011111111111111111011101100010100000000000000000001001111111111111111111111111111111111101000000000000000000000111111101011111111101100111111101101011111111100001111111011001111111110101111111111111111101011111111101100111111101000111111101001011111111101011111111100010111111111111111101111111110101011111111100101111111110000111111101101011010010101011111111111111111101111111110101111111111000011111110100000111100000101111111101100111111111010111111000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111010101010101101010100110010101011111111111111111111111111101010101011010010110010110011111111111111111111111111101010101101001101010010101111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111110010010010110100011111111100100111111101000111111000010100101111111101001011111111111001111111010000000000011111111111111111111111111101111111111111111111111111111111111111111111111101010111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010110000000000000000000100111111111111111111111111111111110000000001000001010100110101111111101011111111111111111010111111111011001111111010010111111111010111111110110011111111101111111111111111111011111111111101011111111100001111111010010111111111010111111110101111111111101111111011111111101011111111101000111110100001011111111101001111111111001111111110101111111111111111110001011010000101111111110000111111101001011111101000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101101001011001010101111111111111111111111111110101010101101010101010100101011111111111111111111111110101011001101010101010010101111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001011010111111111111111110011111111110100111111000000000101111101011101011010111111111110111010000000010111111111011111111110101111111111111111111111111111111111111111111111111111111011111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111110111111111111111111111100000000000000000001010011111111111111111111111110100000000100000000110100110001111111110100111111101100111111111010111111111111111110111111111111010111111111000011111110100101111111110101111111101010111111111111111110111111111010010111111010010111111111000011111110110011111111101011111111101111111111111111111000001111111100011111111010010111111111010011111110110111101000010010000011111111101010111111101100111111101100000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101011101111111111111111111111111110101010110101010011010100101110111111111111111111111111101010101101010101010010101011111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011110010011111110101011111111111011111011111010010100000101111100011100001010001111111111010100000001001111111010101111111110101111111110101111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111110101111111111111111101011010000000100000000000101111111111111111111111010000000001100000100100011101011111111101100111111101000111111101101011111111011001111111110101111111111111111101111111111110011111110110100111111101000111111111101011111111010111010000011111111101111111110110111111110100101111111100101111111110100111111101100111111000010111111111111111010101111111111010111111111000011111010000011010111101010111111111011111110111111111011000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111110101011010101010101010010101011111111111111111111111010101011001011010010101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111000111111110100011111111110101111111101100010010000011111011111110001011011111111010000000000000111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111110101111101011111111111111101010110001010000000001111111111111111111101000000000101000000111000011111111101011111111111111111010111111111101011111111100001111111010001111111111010111111110101111111111111111101011111111101100111111101001011111111100011110000101010111111110101111111111111111101111111111101011111110110101111111101000111110110001001111111011011111111110111110111111111110101111111010000100100010100101111111110000111111101100111111101000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111101010110101001101010100101010101111111111111111111111111110101010110101010101001010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100111110010111111110101011111110110101111111110000010100000001011111111100000111111110111111110000000101111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111110101111111111111111101011111111111111111011101100001010110100111111111111111110110000000010100001001111000011111110100101111111110101111111111010111111111111111010111111111010101111111011010011111110100011111110110101111111101011111111111111111111111111111011011111000100001111111110010111111111000011111110101011111111111111111011111111101010111111101100010011111100001111111010001111111111001111111110101111000101110101101011111111101101111111101001011111111000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101010101010100101010111111111111111111111111111110101010110011010010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010011010011001110101111111111111111111011111111101000000001001100111111111100000101111100011111101000000111111111111111111111001111111110101111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111110101111111111111111101011111010111111111111111011000100111111111111111111111010000000011011000000111010001111111111110011111111110000111111101000111111101101011111111010111111111111111110101111111110110111111111100101111111100000111111101000111111111010111111111011000100111111111110101111111111010111111110100011111110100101111111101101111111111011111010100000111010111111111011001111111010010111111111000110100101000000111111101011111111111111111011111111111011010000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101001010101111111111111111111111111110110011010101010100101010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111001010011111000011111110100011111111101011101000000001111011111111111010110001111011001111101000001111111111111111111110111111111110101111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111101101111111111111111011011111111111111110111010110011111111111111111100000101101100001011111101011110101111111111111111111011111111101100111111111001011111111100011111111011001111111110101111111111111111111111111111101011111111101000111111101001011111111100000101111011011110111111111111101111111110101011111111110101111111100100111111101000111111101000000011111110111110111111111111101111111111010011110000000001011110110101111111110100111111111011111111101100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111111111111111111111111010110101010101010101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011110111010001110101111111110110011111110100001101000000000111111101100111111101000111011111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111101011111110111111111111111110110111111111111111110000001011111111110000010110110101111111101101111111000011111110110101111111101011111111111111111111111111111010111111111010010111111110000111111110100011111110101011111111111111111011111011111010111111111100000101111010001111111010010111111110110111111111101111111111111111101011111111101100111111101000000001001100011111111011001111111110101111111111101000001100011111110101111110110100111111101001011111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111010101101000100010101001010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111010001111111111101111101111111111101110100000010101111111101000111111101000011111111011001100010111111111111110111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101010111111111111111011011111111111111110101011111111111111111010010100111011000001011110101111111111110101111110101011111110100101111111110001111111101000111111111101111111111110111110111111111110101111111111010011111110100101111111110001111111101100111111111011111110100001111010101111111111010111111110010011111110100011111111110011111111101011111011111111111010101100000001001111111010001111111010010111111111000000011010010011111111111111111011111111101100111111101101010000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111010110101000101010101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011001111111100010111111111010011111110110011111011000101111111111111111010111111111100010111111100011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111010111111101111111111111111101100111111111110101010000000010101111111111111111110110010101111111111111111111111111111101101111111101000111111101001011111111101001111111111011111111111111111101111111111110011111111110101111111101000111111101001011110110001011111111110111111111111111110101111111110110011111110100101111111110001111111101101111111111100000000010111111010111111111111001111111111000100001111000011111111110101111111101011111111111111111010111010000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010000010101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011110111111111100001111111111010111111110100011101100000001111111101101111111111011101011000011111110111010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111101011111111111111111110110101001011011111111111111111010111000011111110100011111111101011111111111111111011111111111010111111111101011111111010010111111011010111111110101111111111111111111111111111101001111111101101011111100000011111111010001111111111001111111110101111111111111111101111111111110101111111110000111111101001011100000001011111111010111111111111111110111110000111000011111110110101111111110000111111101000111111111010000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111011000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001001111111011011101011110111111111111111110101110110001010011111111110100111111101000101010100000111111111010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111010111111111111111011001111111111111111010100001111111111111111001110101111111111010011111110100100111111110100111111101010111111111111111110111111111010111111111110010111111111000011111110100101111111110011101101111011111111111111110001011111111011001111111010010111111111010011111110110011111111101111111111111111111011111111111101011110110000010011111100001111111011010111111111000010100011111111101111111111101011111111101100111111101000001100000000010111111111111111111111111111111111111111111111111111111111111111111111111111101000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001101011111111010001001011010010111111110110111111010000011111111111111101011111111101100101011000000011111111010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111101011111111111111111110111111101111111111101000001111111111111100001111111111101111111111111111100011111111110101111111110000111111101000111111111011011111111110111111111111111110101111111110110011111111110001111101110000111111111100110000111010111111111111111110111111111111010111111110100111111110100101111111110101111111101011111111111111111010000000111011001111111110010111111111000101110101000011111111101011111111111111111011111111111010111111000000000100111111111111111111111111111111111111111111111111111111111111111111111110110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001011111111111111010101000111010101111111110010011101000000011111110110011111111101011111111110000010001001111111010010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111011001111111111111110110011111111111011010011111111111000010111111011010111111110110111110111101111111011111111101011111111101100111111111100011111111101001111111111001111111111101111111111111111101011111101101100111111101001001001011101001111111011001111111110111111111111111110111111111110110011111111100101111111101000111111101101011110110000010011111110111111111111111111000100101001000011111110100101111111110100111111111101111111111011101000000000010111111111111111111111111111111111111111111111111111111111111111111110100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000111111111011011111101101011111111111111111101110100100110011111110100101111111110001111110100000010100010011111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111101100111111111111111010101111101111111111111111111010111010110011111111110100101111111111010111111111000011010110110101111111101011111111111011111111111111111010111111111010001111111010010111111111010011111110110011111111101100111111111111111011101001001101011111111100001111111010010111111111010111111110101111111111111111111011111111101101111111101000111111101000000000111011001111111010101111101001010100111111111111110011111111110101111111110000111111101101011011000000000100111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001001100111111101101001111101000001111111011001111111010000011111111111111111011111111101101111011000000001111000000111110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011101101010101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111011111111111011111110101111111111111110110011111111111111101100111101001111111111110011111110111111111111111110101011011110110011111110100100111111110100111111111100111111111011111111111111111110101111111111010011111110100011111111100001111111101100111111101000011111111111111110111111111011001111111110010111111111000011111110110011111111101011111111111111111111111111111011010000010000001111111010010111101000000000111110101111111111101111111011111111111011111111101101001111101000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111010111111110001011111111010010111101000010011111110110011111111101011111111111100000000011110100001011110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011010001000000000000000001010100111111111111111111111111111111101010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111001111111110110111101011111011111111111111111010000100111110110011111010001111111111010111111010001111101111111111101011111111101000111111101001011111111101001111111011011111111110111111111111111111101111111111110100111111110000111111101001011111101101011111111110111111111111111110111111111110110111111110100011111111100101111111101100111111101010111111111100000001011111111011001111111100000100011111000011111110110011111111110011111111101111111111111111111011000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000101111111101100111111111010100101111111111111111110100101010111111111000011111110100101111111110000000000111111110001011111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011000000000000000000000000000000000001001111111111111111111111101010110000000100010100101111111111111111111111111111111111111111111111111010101010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111101011101011111111111100111111111111111011000000010010001111111011010111111011000111111100000011111110110011111111101111111111111111111011111111111101011111111100001111111011010111111111010011111110101111111100111111101011111111101000011111111101011111111100001111111011001111111110101111111111111111101111111111101101111111110000111111101001011111111100000000001011011111111111111100011011001110101011111110100101111111100101111111101000111111101100111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000010101001111111111111111111111111111111111111111111111111111111111111111111111111111111011000100101101111111101000111111111100000011111101001111111010010111111111111111111111111111101011111111000000000000111111111100001111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000100000001010100101011010101010000010100101010100001010101010010101011111111111111111111111111111110101101000101000100010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111110110101111011111111111011111110101111111110110000000000001011111111111111111110101111101101010011111110100011111110110001111111101100111111111010111111111111111110111111111111010111111111000111111110100011111100110011111111101011111100010111111010111111111011011111111010010111111111010111111111010011111110101011111111111011111111111111101010111111111101001100000000001111111010010010001110010111111111101111111111111111101011111111110100111111101001011111111000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001111010011111111111111111111111111111111111111111111111111111111111111111111111111110100000011111111111011111110111111111100000111111100001111101000010111111111010111111110101111111111101010000000000101111111111011000100101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000000000001010110100000100010101000101010011111111111111111010110100010001000101010101001010111111111110110100010100110000111010110000010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111010111111111111111111001111111111111010000001000000011111111011001111111110110101111111111111101111111111110101111111110000111111101001011111111101011111111010111111111111111110101111111110110011101100100101111111110001111100000100111111111010111111111111111111111111111111001111111111000011111110100011111111110101111111101101111111111011111011111111000000001111111011001010001110010111111111000011111110110011111111101111111111111111111010111111111011010100000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111100000111111111111111111111111111111111111111111111111111111111111111111101100010101000101111111101101111111101010111111010011111111111110100101011111111110010111111110100011111110110000000000010011111111111110100101111101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001000000000000000100000001001111111011101010101010111111111111111111111111111111111111111011010101000101000100010100110000010010111111101101011111111011000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111011111110111111111111111111101101111110100100101101011111111010010111111011000011111110110111111110101111111111111111101011111111101100111111101101001111111100001111111011010111111110101111111111101100111011111111101101111100000001011111101000011111111101001111111010101111111111101111111111111111110011111111100101111111110000111111101000111111101100110000000101111110111111001111000111111110110011111110100011111111100101111111101100111111111010111111111100000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111101100010011111111111111111111111111111111111111111111111111111111111011010001001111110011111111110100111111101000111111010001011111111010000111111110111110111111111110110111111110100001010001000011111111111110110000111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000101000000000100000000010010111111111111111111111111111111111111111111111111111111111111111111111110111110101011010100010100111111111111111010010111111111101000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111110011111111000100111111111111111010111111111110010111111111000011111110100011111111110101111111101011111111111111111010111111111011001111111010010111111110010011111110100101111111101011111111101100010011111111111010111111111100001111111010001111111111010111111110101011111111101111111111111111101011111111101100111111111000011111000000011111111010010111110010101111101111111111101011111111110101111111110000111111101001011111111100010000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111110100101001111111111111111111111111111111111111111111111111110110101010010101111111111111011111011111111101010111101001101011111110000001111111010001111111110101111111111101111000000000001010111111111111111101001001100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111010011111111111010000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111110101111111011111111111111111010010001011111111011011111111010111010001111111110101111111110110011111111110101111111110000111111101100111111111010111111111111111111111111111110110111111110100101111110100101111111110000000111101010111111111011111111111111111011001111111011010111111111000011111110110011111111101011111111101111111011111111111010111110110000000011111010010111100001010111111110110011111111101111111111111111101011111111101100111111111100001011000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111110000000101011111111111111111111111111111111111111010110100010100111110100011111111110101111111101011111111111001011011111111000100111111111011010111111010010011111111010001010100000000010111111111111111111010010010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000001001100000000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111111111100000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111101101111111111111111101001100111111111100011111111010010101011111010111111110101111111111111111101011111111101011111111101001011111111001001111111011001111111110101111111111111110110101111111110011111111110000000011101000111111101101011111111010111111111111111110111111111110110111111110100011111110100101111111110001111111101100111111111011111100000100111111000111110000010111111111010011111110100101111111110101111111101011111111111111111010111110101100000001010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111100100111111101101001001000100111111111111111111111111111010110000010100111111111110101011111110110011111111110001111111110000111111111100010011111111111110111111111110101111111110100001010000000000001111111111111111111011000011000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000001010000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111111011111011011111111000111111111111111011111111111011000000111010010111111111000111111110110011111111101011111111111111111011111111111100111111111100011111111010010111111111010011101100110111111111111111111100010011101100111111111001011111111000001111111010001111111111001111111110111111111111111111101011111111110101111111101000111111101001011111000000001111110010110101111111111110101111111110110011111110110101111111110000111111101100101111111010111011000000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100101010101111111111111111111011111111111111111111111111111111110000111111101111111110110100010001010100110010110101010000010000010111111110101111111111111111101111111111101011111111110000111111110001011111111100001111111011001111111110101110100100110000000100001111111111111111111110110100100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000101010000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000111111111111111010000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111101011111111111111111011011111110000111111101101011111111010111110110001111110111111111110110111111110100011111110100101111111110101111111111010111111111111111110111111111111001111111111010111101101000011111110100101111010000101111111111011111111111111111010111111111011001111111011010111111111010011111110110011111111101111111111111111101011111111111101011111101000000011111100000001111011010111111110101111111111111111101011111111101101111111101000111111111001011111101100000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111110101010111111111111111111111111111111111010101010110011111111111111111110101010101011111111111111111111111111111111101000000101111111101101111011110001010100010000010101010011111011001111111011000111111110100011111111110011111111111010100011111111000100111111111011011111111010001111111111010110110010100000000101011111111111111111111111110000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111110001010000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111011111110111111111111111110100100111111101000111111111100011111010100001111111110101111111111111111101111111111101011111111110001111111110000111111111101011111111011011111111111111111101111110101101111111110110101111111000001111111101000111111111100111111111111111110111111111110101111111111010111111110100011111110110101111111110101111111111011111111111111111010000000111111010101111011010111111111000011111110110011111111101011111111111111111111111111101010111111111100010000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111010101110101111111111111111111111111111101011010100101110111111111111111110110100101111101111111111111111111111111111111111111000000011111111110100111111110001011111101001001111111011111111101111111110111111111110110011111110110101111110110100010111101101001111111111111011111111111110111111111011010010010111000000000000111111111111111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111100010011101100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111010111111111111111111111111010111011001101001111111010010111111111010111111110101011111111111111111111111111111100111111101101011111111100001111111010001111111111010101111111101111111111111010000101111111101100111111101001011111111100011111111011011111111110111111111111111110101111111111110101111111110100111111110000111111101100111110100000001111111101011110111111111111001111111110100011111110100101111111110100111111101010111111111111111111111011000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110101101010010101111111111111111111111111110101011010010111111111111111111101011010011001111111111111111111111111111111111111111111111111100010011111111111011111111111100111111101101011111111101001111111111001111111111101111111111111111101011111111110000001111110001011111101001011111111011011111111110111111111100011010000000000000111111111111111111111111111111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010011110100101111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111110101011111100001111110100111111101010111111101100011110111111111110101111111111010011111111000011111110100011111111101101111111111111111111111111111010111111111010001111111110000011111111000011111110110010000011111011111111111111111010111111111101011111111100001111111010010111111111010111111111101111111111111111101011111111101100111111101101011111101000000011111101001111111110101111111111111111101111111111101011111111110100111111101001011111101101011111111011010100000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111010110100101010111111111111111111111111111110110101001110111111111111111111101011010010101111111111111111111111111111111111111111111111111111111110000010110011111111101111111111111111111010111111111011011111111010001111111011010111111110110111111111101111101001011111000101111111111100111111111100011111111100001111101000010000000000000101111111111111111111111111111110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000101000000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001010111111111111110110001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111110110111101100111111110000111111101001011111110000011111111010111111111111111111111111111110101111111110110101111111100100111111101000111111111100111111111110111111111111111110100011111110110011111110100101000011100101111111101100111111111011111111111111111110111111111011001111111111010011111111000011111110110011111111101011111111111111111011111111111010000001011010001111111010010111111111010011111110110111111111111111111011111111101010111111101101011111111100001111000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111110101011010101001011111111111111111111111111101010110101001011111111111111111010110101001100111111111111111111111111111111111111111111111111111111111111111111000001000101111111110001111111101100111111111011111111111111111110111111111111010111111111000011111110110101110100101000001111111011111111111111111010111111111011001111100000000101010000000011111111111111111111111111111111101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000100000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000101111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111110000111111111111111111111010111110100001011111111100001111111010001111111110101111111111101111111111111111101011111111101000111111101001011111111100011111111011001111110010101111111111111111101011000011110101111111110000111111101001011111111101011111111110111111111111111110101111111110110111111110110101111111110100111111101100111111111010111110110000001010011111111011001111111111000111111110100011111110110101111111101101111111111111111111111111111010111111111100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101010101101010100101011111111111111111111111110101011010100111111111111111111111010110101010011111111111111111111111111111111111111111111111111111111111111111111111111110000010011111111101101111111101000111111101001011111111011011111111110111111111111111110101111111110110011000010100001111111110000111111101100111111111010111111111111010010100100100000000011111111111111111111111111111111111010010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000010000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111110100100110100111111101011111111111010000100111111111010111111111011010111111010010011111111010011111111110011111111111011111111111111111010111111111101001111111010010111100010010111111110110111111111000101111111111111101011111111101100111111111101011111111100001111111011001111111110101111111111111111101111111111110101111111110000111111101001011111101000000001011010111111111111111111111111111110101011111110110101111111110100111111101100111111101100111111111011111011000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111110101011010101010010111111111111111111111111111010101100110010111111111111111111101011010011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011101111111111111011111011111111111100111111111100011111111011010111111111001111111111101111111100010100010111111111101100111111101101011111111101001111111010010111100101000000010011111111111111111111111111111111111110110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111011111010001110110101111111110000111111101000000011111100111111111011111111111111111110101111111111010011111110100101111111110100111111101101111111111011111111111111111010111110100011010111111011000011111111000000111111110101111111111011111111111111111010111111111011001111111010010111111110010111111111010011111110101011111111111111111111111111101100111111111100000000011100001111111010010111111110110111111111101111111111111111101011111111101000111111101001011111111101001111101000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111101010110101010101010011111111111111111111111111101010110101001011111111111111111110101101010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101000101111111101101111111101011111111111011111110111111111011001111111110010011111111000011101100000000111111101011111111111111111011111111111101011111111000001110100100000000010111111111111111111111111111111111111111101101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111111111111111111011111110110000000011101100011111111101001111111011001111111110111111111111111111101011111110110101111111110000111111101001011111111101011111111111010111111111111111101111111110000001011110100101111111110000111111101100111111111010111111111111111110111111111111001111111111010011111110100101111111110101111111101011111111111111111010100000001010101111111011001111111110010011111111000011111110110011111111101011111111111111111011111111111101011111111010000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111010110101010001010100101111111111111111111111111110101101010101001111111111111111101110110101010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000101111111110100111111101000111111111100111111111010111111111111111110111111111110110111110101000101111111100101111111101100111111111010111111111110110000111111010111000000010011111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000011111110110011111111101010010010100011111010111111111101001111111010001111111011010111111110110111111111101111111111101111111011111111111100111111111100001111111010010111111111001111111110101111000100001111111011111111110010111111101101011111101001011111111101001111111010111111111110111111101111111110101011111111110101111111110000111111101000111111101000000110111110111111111111111110101111111110110011111110100011111111110101111111101100111111111011111111111111111110110000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010000010001001010111111111111111111111111101010110101010010111111111111111111101011010100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000101011111111011111111101010111111101101011111111100011111111011001111111110101111111111111100010111111111101101111111110001111111101001011111111101000011111010010110100000010011111111111111111111111111111111111111111111111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000001000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100100011111110110001111111110000001111000000111111111011111111111111111110101111111111010111111111000111111110100101111111110010111111101011111111111111111011111111111010001111111011010111111111000011000101000011111111101011111111111111111011111111111100111111111101001111111010001111111111010111111110101111111111101111101111111111101010111111101101011111111000000101111101001111111011001111111110111111111111111111101011111111110101111111110000111111101001011111111101011111101100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0010100101111111111111111111111111110101011010101001011111111111111111110101011010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000100111111101011111111111111111011111111111010111111111010001111111110010111111110100001011110101011111111111011111111111111101010111111111100000011111100001110100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111101111111111100000111110000000111111101001011111111101011111111110111111111111111110101111111110110011111110110101111111110000111111101101011111111010111010001110111110101111111111010011000010100101111110100101111111110100111111111010111111111111111110111111111011011111111011010111111111000011111110110011111110110011111111111011111111111111111011000001011101001111111010010111111111000111111110110111111111101011111111111111111011111111101100111111111101011111111010000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101111111111111111111111111010110101010100101111111111111111111010101101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000001010010110100111111101000111111111010111111111110111110111111111110101111111110000101111110100101111111110101111111101011111111111111111010001111111100011110100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010000111111110110011111111101011000011111100010011111111111100101111111101001111111010001111111011010111111110101111111111111111101011111111101101111111101001011111111000011011011011001111111110101111111110000111100101111111110011111111110100111111110000111111111001011111111010111111111110111111111111111110101111111110100011111111100101111111110100111111101100111110100001001110111111111010111111111111001111111111000011111110100101111111110101111111101011111111111111111010111111111011010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111101011010101010010111111111111111111101011010101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000000000000101111111101000111111101001011111111101011111111010101111111111101100010111111110101011111110110101111111110000111111101000111100001010101001011111000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001010011111111000011111110110000001111111100001111101011111111111111111010111111111011001111111110010111111111000111111110110101111111101011111111111011111111111111111011011101011010001111111010010111111010010011101001001011111111101111111011111111111101111111101101011111111100001111111010001111111011001111111110111111111111111111101011111111110100111111101000111111110000010111111011011111111110101111111111111111101111111110110011111110110100111111110000111111101100111111111010111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111010110101010101001011111111111111111110101101010100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000001010010111111111111111010111111111101011111101100001111111011000001011110110111111111101111111111111111101010111111101100101101011000000000111010000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101000000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010101011111111101111111110100001011111111000011111101000111111111100111111111010111111111111111110111111111110110111111110100011111111100101111111101100111111101010111111111101011110111111111111001111111010000111111100000011111110110101111111101011111111111011111111111111111010111111111011001111111011010111111111010011111110110011111111101011111111111111101011111111111100000101111100001111111010001111111111010111111110101111111111111111101011111111101010111111101001011111111100011111111011000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111011010100010101001111111111111111101110110101010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000010100101101111011111010111011001101000101011111111010000101111111000111111110100011111111110011111111111011111111101000111011000101111010000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000111111011010111111110101011000100111111101001011111101100111111101001011111111100011111111011001111111110101111111110111111101111111111110011111111110000111111101001011111111001001111111010101111111110111100010111101100000111111110100101111111110001111111101000111111101100111111111010111110111111111110101111111111010111111110100011111110100101111111110101111111111010111111000100111110111111111011001111111011010111111111000011111110110011111111101011111111111111111011111111111100111111111010110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101010100111111111111111110101011010101010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100000000000000000000010100000100000000000000001111111110101100010111111110101111111110110011111110110101111111110100111111110000111110100101111110100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111111000111111110100000010111111111110000101011111111111111111011111111111011011111111100001111111010010111111111010111111110101011111111101111111111111111101010111111101001011111111010001111111011000100001111000100010011101111111111111111101011111111110100111111101101011111111101001111111011011111111010101111111111111110101111111110110101111111110100111111101000111110100001011111111010111111111111111110111111111110110111111110100011111110110001111111110100111111111100111111111011111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1001010111111111111111111101101000101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110101100000000000000000000000000000001010001001111111101000001011111001111111110111111111111111111101011111111101100111110100000111110100001011110100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111110111110111111111111000000111111111111110001100100111111101100111111111100111111111110111111111111111111001111111111010011111110100011111110110101111111101101111111111011110100111111111010101111111011000000001111000001000100100011111110110011111111101011111011111111111010111111111101011111111100001111111011010111111111010111111111101111111111111111101011111111101100111111110000011111111100001111111011001111111111001111111111111111111111111111101011111111110100111111101000111111111101011111111011000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111010110100010101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101010111111111111111111111111111111111111111111111111111111111110110001000001001100111111111010111111111010000011111011010111111111010011111110101011111111101111111111111111010010111111000101011110110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111010001111111110110010000011111111111110110101101011111111110100111111101001011111111101001111111011011111111111111111101111111110110011111111110101111111110000111111101001000011111100111111111110111110101000011110110000100000010011111110100101111111110100111111101100111111111011111111111111111110111111111011001111111111010011111111000011111110110011111111101011111111111111101000010111111011011111111010001111111010010111111111010011111110101011111111111111111011111111101010111111101101011111111010100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111011010100010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010101111111111111111111111111111111111111111111111111111111111111110100101110000111111101100111111111111111010000111111110101111111111010111111110100011111110110101111111101100001011111011000011111110100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111111010001111111011000001011111111111111110100101111111101111111011111111111010111111101101011111111100001111111010010111111110101011111111111111101111111111101011111111101101010011111001011111111100001111110000001111111100010000001111111111101111111111110101111111110000111111101001011111111101011111111010111111111111111110101111111110110011111110100101111111100101111111101000111010000100111111111111111110111111111110101111111111010011111110100011111010110101111111101011111111111111111111111111111011110001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101101000101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110010101011111111111111111111111111111111111111111111111111111111111111111011001111101101111111101000111111111001011100001011001111111110111111111111111110111111111111110011111111110000001111101000010111111101000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111111111010000100111111111111111111000101111111110101111111101011111111111111111111111111111010101111111011010111111110000111111110100011111111110011111111101111111111000111111010111111111011001111110000010111111010000000001110110011111111101111111111111111111011111111101100111111111101011111111100001111111011001111111110101111111111111111111111111111101101111111110100111010000001011111111101001111111011011111111110111111101111111110101011111010110101111111110000111111101000111111111100111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110010101111111111111111111111111111111111111111111111111111111111111111111111111011001011111111111111111011111111101101010000011100001111111010010111111110111111111111101111111111111111101001001111101100010111101000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111100011111111010110000010111111111111111111010000111111110110101111111110000111111101001011111111010101111111110111111111111111110111111111110110011111110110001111111110000111111000100111111111011111011111110100000101111111111000010010011000011111110100011111111110101111111111011111111111111111010111111111010101111111010010111111111010011111110100011111111101011111111111111111011111111000001011111111101011111111010001111111010010111111110110111111111101100111111111111101011111111101100111111101101001111111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101100101111111111111111111111111111111111111111111111111111111111111111111111111111110100110101111111101101111111111011111111100000111111111111111111001111111011101011111111000011111110110011111101001011111100001111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111101001111111100000000111111111111111111111010010111101111111111111111101011111111101100111111101001011111111101001111111011001111111111101111101111111111101011111111101101111010010001011111111001011111111100000101111110101111000111000101101111111110110011111110100101111111110000111111101100111111111010111111111111111110111111111111001111111111010011111110100101111111110100111111101010100001011011111111111111111010101111111011001111111110010111111110100000111110101011111111101111111011111111111010111111111010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110010111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111110011111111110001111111101001011111000001011111111010111111111111111111101111111110101011111110100101101001000100111100010100111111000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011011111111111111101100010011111111111111111111111101001110110101111111110011111111111011111111111111111010111111111011001111111010010111111011010111111110110011111111101011111111111101001011111111101011011111111100000111111010001110100100000000111110101111111111111111111011111111101101111111101000111111101101011111111011001111111110101111111111111111101111111110101011111111110101111111110000110000010001011111111011011111111110111111101111111110101111111110100000111110100101111111110001111111101101111111111011111011000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111111111111111111111111111101101111111000001011111111100001111111011001111111110101111111111111111111111110100101101111001010000111011010000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111001011111111010000001001111111111111111111111101101011110110011111110110001111111110001111111101100111111111011111110111111111110111111111111010011111111000011111110100101111111110001011111111011111111111111111100010111111011001111110000000001001111000011111110110011111111101011111111111111111110111111111100111111111100001111111010001111111111010011111110101111111111111111111011111111101010111000010100111111111001011111111101001111111111001111111110101111111100011111101111111111110101111111101000111111101101011111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111010110100101111111111111111101010111111111111111111111111111111111111111111111111111111111111111111111100000011111111110101111111101011111111111010001111111111111010111111111010010111111111010111111110110011111110110101111111101001111111111110010100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111101100111110101000010011111111111111111111111111101001001111111111111111101111111111101101111111101000111111111001001111111011011111111110101111111111111111101111111111110011111111110001111111110000111111101101001100010010101111111111110001001100010110110111111110100011111110100101111111110100111111111010111111111110111111111111111011001111111011010111111111000111111110100011111111101101111111101100000011111111111010111111111011001111111010010111111111000111111100010011111111101111111111111111101011111111111101011111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011001010111111111111111010110100101111111111111111101011010011111111111111111111111111111111111111111111111111111111111111111111101101001011111110110101111111110000111111101000001111111010111111111111111111111111111111001111111111010011111110100101111111100100111111101101011010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101011111111111010000001001111111111111111111111111111110000010111111110110011111111101111111111111111111011111111111100111111111100001111111010001111111111010111111110101111111111111111100101111111101100111111111001010000001100001111111010000000111100000111111111111111111111111111110011111111110100111111110000111111101101011111111010111111111111111111111111111110101111111110110011111110110101111111110000000011101100111111111010111111111111111110111111111111010111111010000011111110100101111111110101111111101011111111111110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010110100101111111111101011010100101111111111111111101011010101111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111101011111111101000001111111001011111111101001111111110101111111111101111111111111110110011111111110001111111110001011010000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101000111110110000010111111111111111111111111111111111110001010111111110100011111110100101111111110101111111101011111111111110111111111111111011001111111111010111111111000011111110110100110011101011111111111111111111000001011011011111111010010001011110000101111111000111111110101011111111101111111011111111101010111111111001011111111000001111111010001111111110101111111110101111111111111111101011111111101100000101101001011111111101011111111101001111111110101111111111111010000011111110110011111111110001111111101000111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011001100111111111111101011010101001111111111111111101011001010111111111111111111111111111111111111111111111111111111111111111111111111111110110111111110110011111111101011111111111011101000001111111010111111111101001111111010001111111111010111111110101110110011101110100101111111101101011100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111101100111010000100111111111111111111111111111111111110100011111111111110101111111111110010111111110000111111101001011111111100111111111010111111111111101110101111111110110011111110100101010111110000111111101000111011000001011111111111111111111101011011000001011111010011111110100101111111110101111111101011111111111011111111111111111010111111111010001111111111001011111111010011111110110011111111101011111111000001111011111111111101011111111100001111111010010111111111010010000111101111111111111111101111111111101100111111101000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011001100111111111111101011010010101111111111111111101011001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111110110011111110100101111111110000101100010010111111111110111110111111111010101111111111010111111111000010110110100010110011101011111010111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001011111011000000010111111111111111111111111111111111111111000011111111010111111111101111111111111011101111111111101101111111101001011111111100001111111011001111111110101111111111111111101010010111110011111111110000111100000001011111111101001111111100001111110000001110111111111110101011111110100011111111110000111111101000111111111100111111111011111111111111111111111111111111010111111110100011111110110101111110100000111111101011111111111111111110111111111011001111111011010011000111000011111110110011111111101011111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111110101011010010111111111111101101010100101111111111111111101011010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111101111101111111111101011111110100000101001010000111111111101011111111011011111111110111110111111111110101111010110110011010111110001111101010000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000110100010101111111111111111111111111111111111111111111010111111111000111111111000011111111110011111111101011111111111011111110111111111011011111111010010111111110010011111111010011111100010011111111101111111111101100010100111111111101001111111010010111111100010111111110110111111111101111111011111111101011111111101100111111101001011111111101001111111011011111111110111111111111111110101011111111110101111110100000111111101000111111101101011111111010111111111111111110101110000110110111111110100101111110110001111111101000111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111110101101001010101111111111101101010100101111111111111111101011010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111010111111110101111111111111011000000101001001010111111101101011111111101001111111011001111111110101111111111010011111011010111101011111010101000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000101111111111111111111111111111111111111111111010001111111110111111111110110111111110100101111111110000111111101100111111111010111111111111111110111111111111010111111111000011101000000101111111110001111110110000001111111011111110111111111010010111111010000101111110010011111111010011111111110011111111101011111011111111111010111111111101011111111010011111111110110111111111010111111111101111111111111111110000111111101100111111111001011111111100001111111011001111111111000011111111111111111111111111101011111111110001111111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111110101011010010111111111111101011010101001111111111111111101011010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111011010111111111000011111110110000010001010000001111111011111111111111111010111111111010001111111010010111111111000011111111000011111111101100111010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111101011000000001011111111111111111111111111111111111111111111111101001011010111111110101111111111111111111111111111101101111111110000111111101001011111111100001111111110101111111111111111111111110000101011111111110101111111000000111111101001011111111101011111010010111111000000111110101111111110110011111110100101111111110101111111101100111111111011111111111111111011111111111110101111111111010011111111000011111110110011110001010011111111111011111110111111111011011111111010010111111010000011111111010011111110101011111111101111111111111111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110101101001010111111111111101011010101001111111111111111101010110010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111111111111111111101111111110100001001100000000000111110000111111111100111111111010111111111111111110101111111110010011111111000011111110100000111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000001111111111111111111111111111111111111111111111111111111111111111111111111111110100000010100111111111111111111111111111111111111111111111111101000111010001111111010000111111111010011111110101011111111111111111111111111111100111111111101011111111100001111111110010111111110100011111111101111101111111100000101111111101101011111111100011111000100001111000000001111111110101111101111111111101011111111110101111111110000111111101001011111111101011111111111111111111111111110101111111110110011111110100101110000000001111111101100111111111010111111111110111111111111111111000101111111000111111110100101111110110100111111101010101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110110100101011101111111111101101010100101011111111111111111010101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010101111111111001111111111101110100000101000001000000011101101111111101101011111111101011111111011001111111110101011001111111110010011111111110001011111000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111101010000000101111111111111111111111111111111111111111111111111111110100111111111111111110101111111110100011111110100101111111110001111111101011111111111111111110111111111111001111111011010111111010000011111110100011111111110000010111111011111111111111111010111110100001001111000000010111111110010111111110110011111111101111111111111111111011111111101100111111111100011111111011011111111011001111111110101111111111111111101111101000010010111111101000111111101001011111111101001111111010101111000100111111111111111111110011111111110101111111110000101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111110110101001010111111111111101100000101011111111111111111111010110101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011001111111011010111111111000101000101110001001010000101111111111111111010111111111101011111111010001111111011010101011110110010001111101111101000111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111101010110101000001001011111111111111111111111111111111111111111111111111111111110000011111111010101111111111111111101111111111101011111111110101111111110000111111101001011111111011011111111110111111111111111100001111111110100011111110100001011111110000111111101100111111111011000011111110010100000011111111010111111111000011111110100101111111110101111111101011111111111111111011111111111011011111111010010111111111000111111110100011111111110001011111111111111011111111111010111111111101011111111010010111000000010111111110110111111111111111101111111111111101110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111110110101010010111111111111101101010100101111111111111111111011010100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111110101111111110110100000110100001011010000000111111101100111111111011111111111111111010111111111111001011001111000101001110100011111100110101000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000011111111111111111111111111111111111111111111111111111111110110001010101001111111111111111111111111111111111111111111111111111111111111111000001001111111010010111111111010011111110101111111111111111111011111111101010111111101100111111111001001111111010001111111010110001011110101111111111111010000101111111101100111111101001011111101000000101111100001111000001011111111111111111101111111110110011111111100101111111110000111111101100111111111010111111111111111111101111111111001111111111010011111110100000011111110001111111101101111111111011111110111111111010111110000000010111111111000011111110100011111111110011111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111011010101010010111111111111101011000100101111111111111111111010110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111011001111111110111110111100010111101000001110100000001111110000111111101001011111111101011111111110111111111011011111111010001110110011101100110101000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111101010111011111111111111111111111111111111111111111111111111111111111111111110010111111111111111011111111011010111111111000011111110100101111111101011111111111111111011111111111010111111111011001111111010000101111111000111111110110000010111101011101111111111111011111111111101000101111100001110100000010111111111010111111110101111111111111111111011111111101101111111101001011111101001011111111110101111111111011111111111111111101111111111110001011111110101111111110000111111101101011111111011011111111010000101111111111110101111111110110101111110110001111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111011000001001010111111111111101101010101011011111111111111111111010101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111010001111111110010111101000010011111100010010110000000111101111111111111100111111111101001111111100001111111010010111111010010111111111101100101010100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111011011111111111111111101111111110101111111110110011111110100100111111110000111111101100111111111111111111111111111110000101111111010011111111000001011110110101111111110101111111111011111110100101111010001111110000010111111110010111111111000011111110100011111111101011111111111111111111111111111010101111111010101111111010010111111111010111111110110111101000001111101111111111101011111111101101011111111100011111111010000100111111001111111111101111111111111111101011111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111011010001001011111111111111101011000101001111111111111111111110110010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111110111111111110110111110000010011111010000101110000000101111111101011111111111111111011111111111011011111111010010111111010000011111110100101111110100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111100011111111010001111111110101111111111111111111011111111101011111111101100111111101101011111111000001111111011001010001110111111111111111010000101111111110101111111110000111111110001011111110001011010010010101000000011111111101111111110110111111110100011111110100101111111110100111111101010111111111111111111111111111010101111111110010111111111000011101000000101111111101101111111111011111111111111111010111111111100000101111010010111111111000111111110110011111111101010100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111101011000001001011111111111111101011010101011011111111111111111010110101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111111111111111111111011011101011111111110101111111110100001101111111111000011110000000001011111110000111111111100111111111010111111111111111011001111111010010111111110100000111110100000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001010000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011111111010111111111011001111111010010011111111000111111110110011111111111111111111111111111010111111111100111111111100010100011010010111111111010000010011101111111111111111101111111111111100111111110001011011001100001010000001001111111110101111111110111111101111111111101101111111110000111111101001011111111101011111111011011111111111111111111111111110101011101000010101111111110001111111110000111111111100111111111010111110000101111110101111111111010111111110100011111111110101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111101101000101001111111111111111101011010101001111111111111111111010110101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111111100111101001111111010001111111010000101111110101111000100100011000000001111101010111111101001011111111101011111111011001111001110101010001111111111101100111111010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001001001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111100111111111011111111111111111110101111111110110111111110100011111110100100111111101101111111111010111111111111111010100000111011001111111110000000001111000101111110110101111111101011111111111111110000111010001011011111000000001111111010010111111111010011111110101011111111111111111111111111111101111111111101011111111100001111111010001011111010101111111110110000101111111111101011111111101101111111101001011111111100011010000001001111111110111111111111111110101011111111110100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101011000001001011111111111111101101000101001111111111111111111110110101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011001111111111111111111111111111111100111110111111111011001111111010010011111111000010100001000011110000000011111111111111111111111111111011011111111100001111001010010010010111010011101101001110110010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000101000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011101001011111111100011111111011001111111110111111111111111110101111111111110011111111110000111111101001011111111101011111000100111111111111111010000100111110110111111111110101111111110001111111101101010101111100001111111110100000001111111110110111111111000011111110100011111110110101111111101111111111111011111110111111111010111111111011001111111010010111111111000000111111110011111111101011111111111111111011111111111101011010000000001111111011010111111111010111111111101111111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1000001001111111111111111101011000101001111111111111111111110110100010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001011111111111111111111111111111111101101111111111010111111111111111100010111111110101110100000000101101100000001011111101100111111111010111111111111111111111111010111001111010111010111111000000010110010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111111011111111111011011111111010001111111110010111111111010111111110101111111111111111111011111111101100111111111001001010010100001111111011010000010010101111111111111111101111111111101101111111110001010101101000001111111100010000010010101111111111111111111111111110110111111111110101111111110011111111101000111111111100111111111110111111111111111110101111111111000000111110100101111111110101111111101100111111111010111111111010000000111111111111001111111011010011111110100011111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1001111111111111111101101010001001111111111111111111010110101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111101101111111111100011111111010010100001110101111111111110000000111111010000000010111110000111111101001011111111101011111111011000011111010010111101111101101001110101100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000101001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001010111111111010111111111111111011101111111111001111111111000011111110100011111111110101111111101011111111111111111110101001011011001111111010000001011111000111111110100011111111101011111111111011111011110101111100001111111101001010000000010111111110010111111110101111111111101111101111111111101111111111101100111111101001001111111101001111111011001111111110111110100101111111101111111110110101111111110000111111101001011111111100000101111010111111111111111110101111111110110011101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111101011000001001111111111111111111010110101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100101111111111111111111111111111111111111111110101111111111010111111111011000000011010010111111111000000000110101010100000000100111111111111111101111111101101001111111100000011111011010111111110110000111110110001000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001001001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001001100111111101001011111111101001111111110111111111111111110111111111110110011111110110101111111110000111111101101011110100001011111111110111010000000111110110111111111000011111110100100111111110101111111100000111100011111111110111110000001011111111011010111111111000011111110100011111111110011111111111011111111111111111010111111111101011111111010010111111010010110100101010011111111101111111111111011111011111111111100111111101100000101111100001111111011010111111110101111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111101101000001001111111111111111111010110101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010111111111111111111111111111111111111111111111110101111010111111111011111110110001011110101111111111010000010110100101101100000000001111101101111111111111111111111111111010101101111010000011111111000000111110100001000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000110001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111011111111111100111111111101001111111100001111111111001111111110101111111111111111101111111111101101111111101000111010010001001111111011010000010010101111111110111111111111111110101011111111110001111110110000111101001001011111111101000000111110111111111111111110101111111110100011111110100101111111110100111111101100111111111011111111111111111010111111111111010111000101000011111110100101111111110101111111101011111111111111111000000101111011011111111010001111111111000011111110100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101011000001001011111111111111111010110101010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010011111111111111111111111111111111111111111111111111110101101001011111111101001110100001001111111111111111101010000010101011111111000000000101110000111111101101011111111100111111111100111110100011111111010001011111000001110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100111111111011111111111111111010111111111011001111111010010111111111000011111110100011111111101011111111111011111011101101001101011111111100000000001010010111111111010111111110110111111111101111111111111111100100111001001101011111111000000000001010001111111111001111111110111111111111111111101111111111110101111111110000111111101001011111111101011111111110111111111111000011101111111110110011111110100101111111110000111111101000101000000000111111111110111111111111111111001111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010001001011111111111111111110110100010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110100111111111111111111111111111111111111111111111111111110110011111010111111111101011111000000001111111011010111111010000011111111101110110000000001001011111111101100111111101101011111111100001110100101001111111101001110110100110000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110000111111111100101111111010111111111110111111111111111111010111111110100011111110100101111111110100111110100001011111111011111100000001111111001111111111010111111111010101111110110101111111101101110101101001011111111111111010110000010011001111111010010111111111010011111110110011111111101111111111111111111010111111111101011111111101001111111100001111111010000011111110101111111111111111111011111111101011111111101101001000000000011111111101001111111111011111111110111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1001111111111111111111110110100010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100101111111111111111111111111111111111111111111111111111111111100101111111111011111111111111000010111111111110001111111111000101111110100011111100000000001111111011111111111111111010111111111011001111110000010111111100010110110101010000010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010111111111101101111111101001011111111100001111111011001111111110101111111111111111111111111111101011111111110000111011000000111111111101000000010101011111111110111111111111111110101111111110110101111111100100100011101001011111101100111111111000010011111111111110101111111111010111111111000011111110100101111111110101111111101011111111111111111010111111111011001111111100010111111111000011111110110011111111101011111111101111111011101000000100111111111101001111111010010111111111010110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111110110100010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101001011111111111111111111111111111111111111111111111111111111111110110011111111101101011111111010010111111010111111111111111110100001111110110011111111000000000011110100111111101100111111111010111111111111101000011111111100010110110010000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000011111101011111111111011111111111111111100111111111100001111111010010111111111010011111110101011111111101111111011101101011100111111111000000001001100001111111010010111111111010111111111101111101111111111101010100011110000111111101001011111111000000101111011001111111110111111111111111111101011111111110011111111110001111111110000111111111100111111111010111111111110111100001111111110110111111110100011111110100101111111110100111111110000000011111011111111111111111110101111111111010010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110101100010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010011111111111111111111111111111111111111111111111111111111111111111110100011111111101100111111111100000111111011001111111011001110110001001111111111111111110000000000110100111111101000111111101101011111111011011101011110101101011110110101010100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111110100101111111101000111111101010111111111111111111111111111111001111111111000111111110100011111110110101111110100001111111111111101000000101111011011111111011001111111011000111111111000011111110110011111110100101110000111111111010111111111100000001111100001111111010010111111011010111111111101111111111111111101111111111101100111111101001011111111100011111111011010000001110101111111111111111101111111111101011111111110001111111100000000011101101001111111011011111111110111111101011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111110100000100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010010111111111111111111111111111111111111111111111111111111111111111111111110110111111011111111111111111100010111111011001111111011010111110000000111111110110011111010000000011011111111111010111111111100101111111100001010001010010101011111010011011010000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101111111101101111111110100111111101001011111111101001111111010101111111111111110111111111110110111111111100101111010000001111111101001000001001100111111111011111111111111111110101111111111010011111110100101111110100100110001101100111111111011111111000000111110111111111011001111111111010111111111000011111110110011111111101011111111111111111011111111111100111111111100000001011010010111111111000111111110110111111111101111111111111110100000000011111101011111111100001111111010010111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1101101010100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001100111111111111111111111111111111111111111111111111111111111111111111111111111110110111110000111111101100111100001010111110111111111110101111110000010111111111000011111111000000010011110101111111111011111111111111111110111110100101001011011010000011011010000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000111110011111111111111111011111111111100111111111101011111111100001111111011010111111110110111111111101111111111110100101010111111101000000101101001011111111100001111111011001111111110101111111111111111101111111111000101100101110000111111101000111110100001011111111010111111111111111110101111111110110011111110100101111111100001111111101100111111111100111111111111111110100001011111001111111111010111111111000011111110110101111111110101000000000011111011111111111010111111111011001111111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101001111111111111111111111111111111111111111111111111111111111111111111111111111111110100111101101111111101000101000001101011111111011001111111110110000000111111111101111111111110000000101110101111111101000111111111101011111111011000001111011001110110011001010000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101011110100011111111100101111111101010111111111111111010111111111010101111111011010111111110010111111111000011111111000101111111111010110000010111111010111111111101001111111010001111111011010011111111010011111111101111010110100101111011111111101100111111110000001111111100001111111011001111111110101111111111111111101111111111101011111111110000111111101001011111101101001110100001011111111111111111101111111110101011111111110101111111110000000000000000111111111100111111111110111110111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101111111111111111101011001011111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111111111111111011101000000001011111111100011111111010000000000011010111111110101111111100000000111011111111101100111111101101011111111100010001011100001110110011010111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111110101011111111110101111111110000111111101000111111111100111111111111111111111111111110101111111110110011101100000101111111110000000000101100111111111011111111111111111110101111111111010111111111000111111110100101010110100001111111101011111111111111110000001111111011011111111010010111111010010011111110110011111111101011111111111111111011111111101010111111111101011111000000001111111010010111111111001111111111101111101111111111101100000000000000111111101001011111111100001111111011000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001010111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101111111110101111111110000000101111111111110111111111111001100000101010011111110100011111111000000001111101011111111111111111011111111111011011011001010010110110010010010000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100101011111111111111111111111111101011111111101100111111111001011111111100001111111011001111111110111111101110110101101011111110100000010111110000111111101101001111111101011111111110111111111111111111101111111110110011001111000100111111110001111111101000110000000010111111111111111111111111111110110111111111000011111110100101111110110100111111101011111111111111111010111010000100101111111011001111111111000011111111000011111111110011111010000000010111111111111010111111111101011111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110010111111111111111011010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101111111110000111111110001010000111101011111111010111111111100010011101111111110101011111110100000010011110001111111101100111111111010111111111111001011001111110010010111000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010011000011111110100011111111101011111111111011111111111111111010111111111011011111111010010111111111000111111100000011111111101011000100111111111011111111111101011111111100001111111010010111111111010111111110101111111010001111000101111111101101111111101001010000000001011111111101001111111010101111111111111110111111111110110111111110110101111111110000111111101001011111111100010111111110111111111111111110101111111110110011111110100101111100000000001111101100111111111011111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010100101111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111110110001001000111001011111111100001111111010010111111110101111111111111111101100000101101101111111101000111111101001011111111101001111010011010010110011000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001110101111111110110010111110100101111111110100111111101100111111111011111111111111111110111111111111010111110101000011111110100000010111110101111111101011111011111111111111111111111011001111111010010111111111000011111010000100000111101011111111111111111111101000000001011111111100011111111010001111111011010111111110101111111111101111101111111111101011111111101100111111101000010111111101001111111011001111111111101111111111111111101011111100000000001111110000111111101101011111111101011110100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011001111111111111110101101001111111111111111111111111111111111111111111111111011001111111111111111111111111111111111111111111111111110110100110101111111101011100001111001011110111111111011011111111010000111111110010011111110100011111100000001011111111111111011111111111100111111111101011111010100000010110010000000000101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111111101111111111111111111011111111110100111111101000111111111001011111111011001111111110111111111011010110101111111010000100111111100101111111101000111111101101011111111010111111111111111111101111111110110111111100000000010010100101111111110100111111101000000101111111111111111111111010101111111011010111111111000111111110110011111110101010111111111011111011111111101000011111111010011111111011010111111011010011111110110011111111101000010001011111111011111111111101011111101100001111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111101011001111111111111111111011010011111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111110100110101111111110001010000101000011111111010111111111111111111000101111110101111111111010011111111000000001111110001111111101010111111111111111110111110100100110100110101000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001010111111111010011111110110011111111101111111111111111101011111111101010111111101100001111111010010111101100010111111110110000010111111111111011111111101100111111101001011111111100011111111010001111111110101111111111111100011100010111110011111111110001111111110000000000111001011111111010111111111110111111101111111110101011111110100011111110100101111111110001111111101100110001011010111111111111111110111111111111010111111111000011111110100001001000010101111111101011111111111111111110111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111101011010011111111111111111011010010111111111111111111111111111111111111111111111110101101001111111111111111111111111111111111111111111111111111111111110001111111111111101010100000101000011111101001011111111101001110110000101111111110111111111111111110100000000111110101111111110000111111111001011111111010000101110101000011000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111101111111111010011111110100011111110110101111111110101111111111011111111111111111110111111111011001111101010010010110000000000111110110011111111101011111111111111111111111111111011011111111010001111111010010111111111000000111100000111111111111111111111111111101000000001001101011111111100001111111010001111111110101111111111101111111111111111101011111111110101111111101000000000101001011111111011001111111110111111111111111111101111111111100001001000000100111111110000111111111101011111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111011010100111111111111111011010100111111111111111111111111111111111111111111111111101011001011111111111111111111111111111111111111111111111111111111111111101100111111101011111110100100111010010111111010111111111101001111110000001111111111010111111110101111101000000101111011111111101011111111101100111111111100010101101000000110100000010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010111111110111111111111111110101111111111110101111111110000111111101000111111101100111111111010111111111111111110101100000000010111111110100101111110110001111111101000111111111010111111111111111011111111111110101111111111000001101100000101111110100011111111101101111000000001001111111111111011011111111011001111111010010011111111010011111110110011111111101111111111111111101100000000111100101111111100011111111010010111111111010111111110101111100000110000111011111111101101111111101001011111111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111010100101111111111111110101101011111111111111111111111111111111111111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111101001011110100101111110100001111110010100111111111110111111111111101000001111111011010111111111000011111010000000111111101011111111111011111111111111111010101000101000000110100000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011111111010010111111111010111111110101111111111111111101111111111101100111111111001011111111100011111111010001110110000000000111111111111111111111111101101111111110100111111101001011111111101001111111010101111111111111111110101101001001011111111110101111111100100111100010000001111111100111111111110111111101111111110101111111111010111111110100011111110100101111111110101111010000000111111111111111011111111111011001111111011010011111111000110100101000001111111101011111111111111111111111111101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111110110101001111111111111111101101001011111111111111111111111111111111111111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111101011111101011111110110000111111000000111111101101011111111011011101001110111111111111111111101111111110000000011111100000111111110100111111111100111111101001001101010100100100000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000111111111111001111111111010011111110100011111110110011111111101011111111111111111011111111111011011111111100001011000000000101001111010011111111101011111111111111111011111111111100111111111100011111111100001111111011010111110100100001011111101111111111111111101011111000010000001111101001011111111101011111111011011111111110111111111111111110101011111111110101111111110001111100000001011111111100111111111010111111111111111110101111111110110011000010100001111111100100111111101100111111111010110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110110101001011111111111111101101010010111111111111111111111111111111111111111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111101110100101111110100000111111111101011111111100001110000101001111111111001111111110111111100000010111101011111111101100111111101001011111111100001100110000000101000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111110111111111111111110111111111110110011111110100101111111110001111111101000111111111010111111111011111110110000000100000100111111000111111110100101111111110100111111101010111111111011111111111111111010101111111010001110110101000000111111010011111110110011111111101100001100010011111010111111111101001111111100001111111010010111111111010111111111101111111111111111101011101000000001111111101001011111111100001111111011010111111110101111111110000011100101111111101101111111110000111111101000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111101101010010111111111111111011010100111111111111111111111111111111111111111111111111111101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111011010011111110110101000001110101100000111011111111111111111010111111000000001111111011000111111111000011110000000011111111101111111111111111111010111111101100010101010000000101000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000101111111111111111111111111111111111111111111111111111111111111111111111111111111111010010111111010001111111011001111111110101111111111101111111011111111101101111111101000111111101001011111111101001110100000010011010011101111111111111110110111111110110101111111110000111111101100111111101010111111111110111111111110110111000101111110100011111110100101111111100000011010000100111111111011111111111111111110101111111111001111111111000111111111000011111111110101111111110000000011111011111110111111111011011111111010001111111010010011111010000110100101110011111111101111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111101101000100111111111111111111010101011111111111111111111111111111111111111111111111111010110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111110110101000100110100101001010000111111101011011111111111000000111111111110111111111110110011111100000001111111110101111111101101111111111011111111000000110101000101000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111101000011111111011011111111010010111111111000111111110110011111111101011111111111011111011111111111100111111111100001100000000010101011111010111111110101011111111101111111011111111101011111111101000111111111001001111111101001111111011010111000101101111111111111111101011111111110001011010000000111111101001011111111101011111111010111111111111111110101111111110110011111110100101111110100000000111101100111111111010111111111111111110111111111110101111111100000011000110100011111111110101111111101011111010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111011000100111111111111111110110101001011111111111111111111111111111111111111111111111110101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111101111111111000100101011101000000100111111111001011111111100010001011011001111111110101111111111111010000000111111110101111111110001111111101000111110100001010101110000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111110100100111010111111111110111110111111111111001111111111010011111110100101111111110101111111101011111111111011111100000000001011000101111010010111111111000011111110110101111111110011111111101011111111111111111010111111111011001111111010010111000010010111111110110111111111101111111100011011000100111111101100111111111101011111111100001111111011001111111110101111111111101111111111111110000000001111101000111111101001011111111100011111111011011111111111101000001110010110101011111110110101111111110000111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111011000001001111111111111110101101010011111111111111111111111111111111111111111111111111101101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100011000011111111000101111111101100000111111111111010111111111011011100001010001111111010010111111111010011000000001011111111111111111011111111101100111111110000010000100000010100000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111110000011111001011111111101001111111111011111111111101111101111111110101011111111100101111111110000111111101101001100000001011111010010111111111111111110110111111110110011111110100101111111101100111111101100111111111011111110111111111010001010010111010111111111000011111110100101111100010100000101111011111111111111111010111111111011011111111010010111111110010011111110110011111110101100000000010111111011111111111100111111111101001111111010010111111010000001011010000111111110101111111011111111101101110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111011010001001011111111111111101011010010111111111111111111111111111111111111111111111111111011010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010111111111000101111111110000000101101100111111111011111111111010000010101111111110101111111111010010100000000101111111110101111111101011111111111111110001010100110000010100000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001111111111111111111111111111111111111111111111111111111111111111111111111111100010111111010111111111100011111111010010111111111010111111110101111111111111111111011111111101010111111101000000000010000001010001010001111111111001111111111101111101111111111101011111111110100111111101001011111111100011111111011001100111010010111111111111110101111111110110011111100000001000101110000111111101100111111111010111111111110111111101111111110110111111111000011111110100000000000000100111111101101111111111011111110111111111010111111111111000000111010000111111110100011111111110011111110110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111110110000010010111111111111111011010100101111111111111111111111111111111111111111111111111110110101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000111111111111000101111111110101000000110000111111101001011111111100000101111010101111111111111110101111101000000011111110110101111111110000111111101100111001010001000000010010000100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000111111111111111111111111111111111111111111111111111111111111111111111111110001001010111111111111111110111111111010101111111111010111111111000011111110100011111111110011111111111010110000000001001010110000111010011111111010010111111111000111111110110011111111101111111011111111111011111111101101011111111100010001111000010111111111010111111110101111111111101000001010100101110101111111101001011111101001011111111101001111111110101111111110111111101111111110110000000001010101111111110000111111101101011111111010111111111110111110100101111000010111111110100011111110100101111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111110000010101111111111111111111010001001111111111111111111111111111111111111111111111111111101101010011111111111110101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101011110110010100100101111111110110000001011111111101010111111111100010001011010001111111011001111111110110000000011111111101111111111101101111111101000111010010000010101010100000100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000111111111111111111111111111111111111111111111111111111111111111111111111000101101000111111101001011111111011011111111110111110101111111110101111111110110011111110110001111111110000000101010001011111100101111111111111111110101111111111010111111110100101111110110101111111101100111111111010111111111111111010110011110001001111111010010011111111000011111110110001011110100001111111111111111011111111111011011111111101001111111010010111111111010111111110101110100000000000111011111111101011111111101101011111111000001111111100001111000011010001011110111111111111111111101011111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111110101100010100111111111111111110110001010011111111111111111111111111111111111111111111111111111011010010111111111111101011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111000010100100100101111111110000000011111011111111111011111011101100010011001111111010010111111111000000000100110011111111101011111111111111111110111010010000000000010100000000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000111111111111111111111111111111111111111111111111111111111111111111111010010111101010111111111101011111111100001111111011001111111111001111111110111111111111111111101011111110110001001111000001011111000000011111111011001111111110111111111111111110101111111111110101111111110001111111101001011111111101011111110101000000111111111110101111111110110111111011000001011110100001111111110100111111101010111111111111111110111111111011001111111011010011111111000101000001000001111111110011111111101111111111111111111010111111111011001010010010000001011111000011111110110011111111101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111101011000100101111111111111111101100010010111111111111111111111111111111111111111111111111111111010100101111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111101111000100110011111111110000000001010001011111101100111111111100000011111111111111111111111110110111000001000101111110100101111111110100111111111100000000000000010011000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001011111111111111111111111111111111111111111111111111111111111111111101001010011111111111111111011111111111010111111111011001111111010010111111111000011111110110011111111101011010111111010000101111011001100111111111100001111111010010111111111010111111110101111111111111111101011111111101100111111101001011110110000000101111011001111111110101111111111111111110000111110100000111111110001111111101001011111101101011111111011011111111111111110111111111110110010000100000011111111110001111111110000111111101100111111111010111110111100001110100001111111010111111110100011111110100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111011000001001011111111111111101011000100111111111111111111111111111111111111111111111111111111110101001011111111111111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000111111110100101111111111111101111000000000101111111101000111111111100000100111010011111111110101111111111000001011111111111101011111111110101111111110000000000000000010111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111110100001110000111111101000111111111100111111111110111111111111111110101111111111010111111111000011111110100001111111101000001111101001011110111111111011111111111011001111111111000111111110100011111110110101111111101011111111111111111111111110101100000011111010010111111010010111111111000111111001010011110001011111111111111111101010111111111001011111111100001111111010001111111110110111111000010010000011111111101011111111101100111111101001011111111101011111111100001110100000101111111111111110101111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010000001011111111111111111011010001011111111111111111111111111111111111111111111111111111111101010011111111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000101111111000000111110110011111111110000000000111111111111111111111011010001011010001111111010010111111111000001011111101111111111111111111111111111111010101101000000010111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001011111111111111111111111111111111111111111111111111111111111111010010111101011111111101100111111101001011111111101001111111011001011111110111111111111111111101011111111110011111111100001011111110000111111111101011111111010111111111111111110101111111110110011111110100101111111110000111111101100111111111101011010010111111110111111111110101111111111010111101000000011110000000101111111101011111111111011111111111111111010111111111011010111111010010111101000000000010110110011111111101111111111111111111011111111111101011111101000001110100000010111111111010111111111101100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010011111111111111111110110001001111111111111111111111111111111111111111111111111111111011010100111111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111110100001111110100101111110100001000000010000111111111100111111111100010011111111111110101111111011000000010111000011111110110101111111101101111111101110110000010111000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111101001001011111111111011111111111111111011111111111101011111111100000111111010010111111111010111111111101111111111111110110000111111000100111111101101011111111100001111111011001111111110101111111111111111111111111111101011111111101000111111101001011000001100011111111010101111111110111111101111101001010111110001010101111111110001111111101000111111111100111111111110111111111111111110101110100001000000001110100011111110110101111111101101111111111011111111111110100100111111000011001111111111010011111111000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111110110100010011111111111111111111111111111111111111111111111111111110110101001111111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001110110000111111111111111111101011101100000001001111101001011111111100000101111010101111111111111111101000010111101011111111110101111110110001111111101000110000000100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011111111111111111111111111111111111111111111111111111111110100100110101111111110100111111101100111111111011111111111111111011001111111011001111111111010011111110100011111110110100100011101010001111111111111010111111111011001111111010010111111110010111111111010011111111101011111111111011111111111111111100101000111101001111111100001111111011010111111110100000111110110001001111111111101011111111101100111111101001011111111101001111111011011111111111000101110000001111101011111111110010111111110000111111101000111111111100000101111010010111111111111110101111111111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111101101000101111111111111111111111111111111111111111111111111111111101100010111111111111111101101001111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010111110000010111111110101011111111111110110000000101001100111111101101000000111100001111111010010111101100000011111111101111111111111111101111111111101000110000000000000000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011111111111111111111111111111111111111111111111111111111010000011101111111111110101111111101000111111101001011111111101001101011110111111111111111110101111111110110011111110110000000111110000001111101100111111111010111111111111111111111111111110110111111111000011111110100101111111110100111111101101111111110000111111111111111111011111111011010111111110000000111110100001011111110011111111101111111011111111111010111111111101011111111100001111111010000011110000010111111111101111111111111111111011111111101100111111101100000011111100010111111011001111111110101011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111011010101011111111111111111111111111111111111111111111111111111111011010100111111111111111011010011111111111111111111111111111111111111101010101111111111111111111111111111111111111111111111111111111111111111111111111111111010111110101111110000010111111110100011111110100101111011000000000001001011111111101100010010111111111011010011011010000101111110100011111111110011111111101011111111110000000101000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011111111111111111111111111111111111111111111111111111101001001111111111101011111111111111111011111111111100111111111100010011111100001111111011001111111110101111111111101111101100010111110001011111101000111111101001011111111101001111111110101111111111111111111111111111110011111111110101111111110000111110100001011111111010111111111011111110111111111110100000111111000001011110100101111111110001111111101101111111111010111111111111111110111111111000010111000000010011111110100011111111110101111111101011111111111111111100001111101000011111111010010111111110000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111010001001111111111111111111111111111111111111111111111111111111110110101011011111111111110110100101111111111111111111111111111111111101011001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111110001001111111110101111111111110101111110110001010001000000010100101100000011111110111011010101011111000001111110110011111110100101111111110100111111110000000110100000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001001111111111111111111111111111111111111111111111111111000100111011111110110101111111110101111111101011111111111111111100010111111011001111111010010111111111000111111110110011111000000111110001111011111011111111111100111111111100011111111010010111111111010111111110110111111111101111111011111111101010111110000101011111101100011111111100001111111111001111110001011111110001011111101111111111110101111111110000111111101001011111111101011111111010110001011111000001101111111110110011111110100101111111110000111111101000111001001010101000111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0110100010111111111111111111111111111111111111111111111111111111111110100001111111111111111110101001111111111111111111111111111111111111110101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111111010000001011111001111111111101111111111111111101011111110101101000100000000000001010100010101001011001111000001001111111111111111101111111111110101111111110000000010100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111101010111111111111110110011111111110101111111110000111111101101010100111010111111111111111111111111111111001111111111000011101000000100100011110101111111101010111111111110111111111111111111011111111011010111111111000011111110110101111111101101111111111100001011111111111010111111111011001111111010010111110000010011110000010011111111101111111111111111111011111111101100111111101100001111111100000001111010000101111110101111111111101111111111111111101011111111101000110100111000000001111101001111111010101111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1010101111111111111111111111111111111111111111111111111111111111101010101111111111111101011010101111111111111111111111111111111111111101011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111011010100001111000111111110100011111111110011111111101011111111111110111010110100000101001011111010001111100000010111111110110011111111101011111111111111100000000111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111111111111111111111111111111111111111110110101011111111110101111111111111111101011111111101010111111101000010011111001011111111100001111111111011111111110111111111111110001010011000011100101111111110000111111101101011111111011011111111110111111101111111110101111111110110011111110110100111111110001011111111100111111111011111111111111111110101110100101010111101000000011111110100101111111110101111111101011111111111111111011111111111100000011111010000011111110000111111110110011111110101011111111101111111110100101111100000101111100011111111010010100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111011010101011111111111111110110101011111111111111111111111111111111111101011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101111111111010010110101111111110110011111110100101111111110001111111101100111111111010101111111111111110111111110000010011111111010011111110100101111111110101110000000010110000000000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111011000011111111111111000011111110110011111111101011111111111010110001001111111011011111111011001111111010010111111111010111111110100000111010010111111111111111101010111111101001011111111100001111111010001111111111001111111110101111111111111111101011111111110000111111101001011111111001001111111011001111111111010011111111110001001111111111110011111110110001111111110000111111101101011111111010101100001110111100010111111110110111111111000011111110100101111111110100111111000001111111000101111111111111111011000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110110101010111111111111111110101010111111111111111111111111111111111111110110010101111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111010000111111110101111111111111111111011111111101100111111101000111111111001011111111011001111111010101000001111111111101111111110110011111111100100100001000000110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000001111111111111111111111111111111111111111101101011111111111111110110111111110100011111111100001111111110000010011111010111111111011111110111111111010101111111110010111111111000101111100000101111111110011111111111111111111111111111010111111111011010111111010010011111111000111111110110011111111101110100101111111111010111111101101011111111100001111111010000011111011000001011110101111111111111111101111111111101101111111101000111111101000010000111101010000001111001111111111101111111111111111101011111111110100111010000000111100000001011111111011011110100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111101101010010111111111111101101010011111111111111111111111111111111111111101011001011111111111010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111010000011111111010111111110110011111111101011111111111111101011111111111100111111111100011111111010010000001111010111111110101111111111111111111111110001000100101000000000000000000000010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111110100101111111111110101111111111111111101111111111101011111011000000101111110001011111111101011111111010111111111110111111101111111111000101111100000011111111100101111111110000111111111100111111111010111111111111111110101111111111010011111110100101111110100000010011101101111111111011111111111111111010111111111010010111111011000000111111000011111110110011111111101011111111111111111011111111111010000101111100000001011010010111111111010011111110110111111111101111101011111100010101101000010101011111111100001100001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111101011010100111111111111111010110101011111111111111111111111111111111111111011010010111111111110101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111000101111111010111111111000011111111100011111111110101111111101010111111111111111110111111111011001100010011010111111111000011111110100011111110100001000011110000000000000000000100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100010111111111111111111111111111111111111100001111111111111010010111111111010011111110101111101011010001001111111111111101111111111101011111111100001111111010001111111111001011010111110001011111111111101011111111101000111111101001001111111101001111111011001111111110101111111111111111101111111111110000001111110000111111110001011111111101011111111010111110010111111110100000111110110111111110100101111110100100111111101000111111101010111100000011111111000001011111001111111111010111111111000011111110100011111111110000111111110001011011111111111011000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111010110001001111111111111110101101001011111111111111111111111111111111111110110100101111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101001110100001011111111111111111111111111111110011111111110101111111101000111111111101011111111010111111111010010110101111111110110111111110110101111111110001010011110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111110110100111111111111111110101111111111000111111111000101010000000001111111101101111111111011111110111111111011011111111011001111111011000010010111000001111110110011111111101011111111111111111010111111111101011111111010001111111010010111111111010111111111101011101000001111101011111111111100111111101001011111111100001010001010001111100001001111111111111111101111111111101101111111110100111111101001001100001001001110000001010011111110111111101111111111101011111110110011111110100000111111100001011111111100111011000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111110101101010011111111111111101101010011111111111111111111111111111111111111111101010011111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111110000010111111111010011111110110111111111101111101011111111101101111111101101011111111100001111111010010011111110101111111111111111101111111110100101000111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100001111111111111111111111111111111011010011111111111011011111111110111111111011101100000001010010110101111111110100111111101100111111111100111111111010111110111111111111001100010111000101111110100101111110110101111111101100111111111011111111111111111010101111111111010111111111010011111111000011110001010101111111101011111111111111111010111111111011011001011010001110110000010111111111010011111111110111111111101111111011111111101101000000111101011100000000000011111011010111111111001111111111101111111111111010000011111111000100111111101001010100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111101101000100111111111111111011010100111111111111111111111111111111111111111010110100111111111111110100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011111111000010111111111010111111110100011111110110011111111101011111111111011111011111111111100111111111010000111111010010111111111000011111110110110100100100011111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111101101001111111111111010001111111011010101010000000000000000101111111111111111101011111111101100111111101101001111111101001111111011001111111100010111000011111110101111111111110101111111110000111111101001011111101101011111111110111111111111111111101111111110110011000010100101111111110000111111101000111111111010111111101001011010111110100001001111111111000111111110100101111111110100111111101011111010000001011010101000010011001111111011010111111011010011111111000011111110110000001111101010000011111111111010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111011000101011111111111111110110001001111111111111111111111111111111111111110101101001111111111111011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001010111100010011111110101111111110101011111111100101111111110000111111101100111111111010111111111110111111000011111110101111111111010111111110100100100011000101111010000000000000010000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100001111111111111111111111111110100101111111111111111010111011010000000001010000000000000111000011111110110011111111101011111111111111111010111111111101001111111010001111101000010111010010110011111111101111111011111111101011111111101100111111111100011111111100001111111111010111111110101111111010010111111111111111101011111111101000111111101001011111110001011111111011000101111110111111111111111111110111111110110101111111110000101001010001011111110000001111111010111110111111111110101111111110110111111110100001011110110000010111101100111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111110110101001011111111111111110100010111111111111111111111111111111111111111111011010010111111111110110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111000100001111111110101111111111111111111111111111101011111111101000111111101001011111111101001110100001011111111111111111111111111110101111000111000101111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011111111111111111111111111011001010111111111011011111111101010100101110101000000000001110110011111111100101111111110001111111101100111111111010111111111111111110101111101000001010010111000111111111000011111111110101111111101011111111111111111011111111111011001111111010010111111111000011111100000011111111101011111111111011111011111111111010111110110000001111111010000011111011010111111110110111111111101111101111111111101010100100110000111110100000011011111100011111111011001111111110111111111111111110100001111111110000001111110001010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111101100010010111111111111111101000101111111111111111111111111111111111111111110110100101111111111101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011110100000001111111111000111111110100011111111110011111111111111111111111111111010111111111101011110100000001111111010010111111110110111111111000011000111111110100000000000000000000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101001111111111111111111111111111111100111111111101011111111110111111111111110000000000111111111111111111101111111111110101111111110000111111101001011111111101011111111110110001011010010110101111111111110011111110110101111111110000111111101100111111111010111111111111111111111111111110101111110101000011111110100101111111110100111111101010111111111011000101111111111010000011111110001111111111000111111110100011111111110011111110101011010011111011000000111111111101011111111010001111111110010111111111010100000011101011110001011111101000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
);

begin

PROM_OP <= mem(conv_integer(addr)); 


end Behavioral;
